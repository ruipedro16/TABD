<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Federacao Portuguesa De Natacao" version="11.69847">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Vila Nova de Famalicão" name="XXII Campeonato Nacional Masters de Verão - OPEN " name.en="XXII Portuguese Summer Masters Championships - OPEN" course="LCM" deadline="2021-06-25" entrytype="OPEN" number="9" organizer="Federação Portuguesa de Natação" organizer.url="https://fpnatacao.pt/evento.php?codigo=559" result.url="https://fpnatacao.pt/Resultados/provas2021/09cnmastersOPEN/#" startmethod="1" timing="AUTOMATIC" type="POR.MNP" withdrawuntil="2021-06-26" nation="POR" maxentriesathlete="5">
      <AGEDATE value="2021-01-10" type="YEAR" />
      <POOL name="Piscina Municipal de Vila Nova de Famalicão" lanemin="1" lanemax="8" />
      <FACILITY city="Vila Nova de Famalicão" name="Piscina Municipal de Vila Nova de Famalicão" nation="POR" />
      <POINTTABLE pointtableid="1124" name="DSV Master Performance Table" version="2020" />
      <CONTACT city="Cruz Quebrada- Dafundo" email="inscricoes@fpnatacao.pt" name="Eduardo Miranda" phone="+351214158190" street="Moradia do JAMOR" street2="Estrada da Costa" zip="1495-688" />
      <QUALIFY from="2019-01-01" until="2021-07-08" />
      <SESSIONS>
        <SESSION date="2021-07-09" daytime="10:00" endtime="19:59" name="1ª Jornada-1ª sessão" number="1" warmupfrom="08:30" warmupuntil="09:45">
          <EVENTS>
            <EVENT eventid="1060" daytime="10:00" gender="F" number="1" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1076" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43959" />
                    <RANKING order="2" place="2" resultid="43294" />
                    <RANKING order="3" place="3" resultid="42462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1077" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43660" />
                    <RANKING order="2" place="2" resultid="41540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43245" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43525" />
                    <RANKING order="2" place="2" resultid="42695" />
                    <RANKING order="3" place="3" resultid="43397" />
                    <RANKING order="4" place="4" resultid="43043" />
                    <RANKING order="5" place="5" resultid="43333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1080" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43276" />
                    <RANKING order="2" place="2" resultid="43499" />
                    <RANKING order="3" place="3" resultid="42028" />
                    <RANKING order="4" place="4" resultid="41944" />
                    <RANKING order="5" place="5" resultid="43625" />
                    <RANKING order="6" place="6" resultid="43455" />
                    <RANKING order="7" place="7" resultid="43210" />
                    <RANKING order="8" place="8" resultid="43179" />
                    <RANKING order="9" place="-1" resultid="43767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42043" />
                    <RANKING order="2" place="2" resultid="43220" />
                    <RANKING order="3" place="3" resultid="43432" />
                    <RANKING order="4" place="4" resultid="42173" />
                    <RANKING order="5" place="5" resultid="43678" />
                    <RANKING order="6" place="6" resultid="41934" />
                    <RANKING order="7" place="7" resultid="44012" />
                    <RANKING order="8" place="8" resultid="43899" />
                    <RANKING order="9" place="-1" resultid="41960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43327" />
                    <RANKING order="2" place="2" resultid="43875" />
                    <RANKING order="3" place="3" resultid="42689" />
                    <RANKING order="4" place="4" resultid="43122" />
                    <RANKING order="5" place="5" resultid="41755" />
                    <RANKING order="6" place="6" resultid="43234" />
                    <RANKING order="7" place="7" resultid="43649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41743" />
                    <RANKING order="2" place="2" resultid="43288" />
                    <RANKING order="3" place="3" resultid="43643" />
                    <RANKING order="4" place="-1" resultid="43569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="1085" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="1086" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="1087" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="8891" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="14943" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45139" agemax="-1" agemin="-1" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43959" />
                    <RANKING order="2" place="2" resultid="42043" />
                    <RANKING order="3" place="3" resultid="43660" />
                    <RANKING order="4" place="4" resultid="43276" />
                    <RANKING order="5" place="5" resultid="43220" />
                    <RANKING order="6" place="6" resultid="43525" />
                    <RANKING order="7" place="7" resultid="42695" />
                    <RANKING order="8" place="8" resultid="43499" />
                    <RANKING order="9" place="9" resultid="43294" />
                    <RANKING order="10" place="10" resultid="41540" />
                    <RANKING order="11" place="11" resultid="42462" />
                    <RANKING order="12" place="12" resultid="43327" />
                    <RANKING order="13" place="13" resultid="43432" />
                    <RANKING order="14" place="14" resultid="43397" />
                    <RANKING order="15" place="15" resultid="43875" />
                    <RANKING order="16" place="16" resultid="42028" />
                    <RANKING order="17" place="17" resultid="42173" />
                    <RANKING order="18" place="18" resultid="43678" />
                    <RANKING order="19" place="19" resultid="41934" />
                    <RANKING order="20" place="20" resultid="41944" />
                    <RANKING order="21" place="21" resultid="42689" />
                    <RANKING order="22" place="22" resultid="43625" />
                    <RANKING order="23" place="23" resultid="43043" />
                    <RANKING order="24" place="24" resultid="43122" />
                    <RANKING order="25" place="25" resultid="41743" />
                    <RANKING order="26" place="26" resultid="43455" />
                    <RANKING order="27" place="27" resultid="44012" />
                    <RANKING order="28" place="28" resultid="43245" />
                    <RANKING order="29" place="29" resultid="43899" />
                    <RANKING order="30" place="30" resultid="41755" />
                    <RANKING order="31" place="31" resultid="43234" />
                    <RANKING order="32" place="32" resultid="43649" />
                    <RANKING order="33" place="33" resultid="43210" />
                    <RANKING order="34" place="34" resultid="43288" />
                    <RANKING order="35" place="35" resultid="43333" />
                    <RANKING order="36" place="36" resultid="43643" />
                    <RANKING order="37" place="37" resultid="43179" />
                    <RANKING order="38" place="-1" resultid="43569" />
                    <RANKING order="39" place="-1" resultid="43767" />
                    <RANKING order="40" place="-1" resultid="41960" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45074" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45075" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="45076" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="45077" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="45078" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1058" daytime="11:00" gender="M" number="2" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="8892" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42812" />
                    <RANKING order="2" place="2" resultid="41731" />
                    <RANKING order="3" place="3" resultid="43483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8893" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42010" />
                    <RANKING order="2" place="2" resultid="43308" />
                    <RANKING order="3" place="3" resultid="43269" />
                    <RANKING order="4" place="4" resultid="43951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8894" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42467" />
                    <RANKING order="2" place="2" resultid="43789" />
                    <RANKING order="3" place="3" resultid="43816" />
                    <RANKING order="4" place="-1" resultid="41828" />
                    <RANKING order="5" place="-1" resultid="42049" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8895" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42987" />
                    <RANKING order="2" place="2" resultid="42064" />
                    <RANKING order="3" place="3" resultid="43693" />
                    <RANKING order="4" place="4" resultid="41749" />
                    <RANKING order="5" place="-1" resultid="41955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8896" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41965" />
                    <RANKING order="2" place="2" resultid="43597" />
                    <RANKING order="3" place="3" resultid="42955" />
                    <RANKING order="4" place="4" resultid="42093" />
                    <RANKING order="5" place="5" resultid="42427" />
                    <RANKING order="6" place="6" resultid="43376" />
                    <RANKING order="7" place="7" resultid="43417" />
                    <RANKING order="8" place="8" resultid="43988" />
                    <RANKING order="9" place="9" resultid="43722" />
                    <RANKING order="10" place="10" resultid="43324" />
                    <RANKING order="11" place="-1" resultid="43984" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8897" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43319" />
                    <RANKING order="2" place="2" resultid="42179" />
                    <RANKING order="3" place="3" resultid="43761" />
                    <RANKING order="4" place="4" resultid="42706" />
                    <RANKING order="5" place="5" resultid="43350" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8898" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43610" />
                    <RANKING order="2" place="2" resultid="43799" />
                    <RANKING order="3" place="3" resultid="43056" />
                    <RANKING order="4" place="4" resultid="43189" />
                    <RANKING order="5" place="5" resultid="43069" />
                    <RANKING order="6" place="6" resultid="43013" />
                    <RANKING order="7" place="7" resultid="43810" />
                    <RANKING order="8" place="8" resultid="43182" />
                    <RANKING order="9" place="-1" resultid="41534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8899" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42972" />
                    <RANKING order="2" place="2" resultid="41684" />
                    <RANKING order="3" place="3" resultid="43519" />
                    <RANKING order="4" place="4" resultid="43488" />
                    <RANKING order="5" place="5" resultid="43880" />
                    <RANKING order="6" place="6" resultid="43451" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8900" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43128" />
                    <RANKING order="2" place="2" resultid="42493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8901" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41658" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8902" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="41652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="8903" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="8904" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="8905" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45138" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43610" />
                    <RANKING order="2" place="2" resultid="42987" />
                    <RANKING order="3" place="3" resultid="42972" />
                    <RANKING order="4" place="4" resultid="42812" />
                    <RANKING order="5" place="5" resultid="42010" />
                    <RANKING order="6" place="6" resultid="41684" />
                    <RANKING order="7" place="7" resultid="43308" />
                    <RANKING order="8" place="8" resultid="43319" />
                    <RANKING order="9" place="9" resultid="41965" />
                    <RANKING order="10" place="10" resultid="43799" />
                    <RANKING order="11" place="11" resultid="43597" />
                    <RANKING order="12" place="12" resultid="43269" />
                    <RANKING order="13" place="13" resultid="41731" />
                    <RANKING order="14" place="14" resultid="42955" />
                    <RANKING order="15" place="15" resultid="42093" />
                    <RANKING order="16" place="16" resultid="42179" />
                    <RANKING order="17" place="17" resultid="42427" />
                    <RANKING order="18" place="18" resultid="42064" />
                    <RANKING order="19" place="19" resultid="43376" />
                    <RANKING order="20" place="20" resultid="43519" />
                    <RANKING order="21" place="21" resultid="43951" />
                    <RANKING order="22" place="22" resultid="42467" />
                    <RANKING order="23" place="23" resultid="41658" />
                    <RANKING order="24" place="24" resultid="43417" />
                    <RANKING order="25" place="25" resultid="43988" />
                    <RANKING order="26" place="26" resultid="43056" />
                    <RANKING order="27" place="27" resultid="43693" />
                    <RANKING order="28" place="28" resultid="43189" />
                    <RANKING order="29" place="29" resultid="43722" />
                    <RANKING order="30" place="30" resultid="43761" />
                    <RANKING order="31" place="31" resultid="43789" />
                    <RANKING order="32" place="32" resultid="42706" />
                    <RANKING order="33" place="33" resultid="41749" />
                    <RANKING order="34" place="34" resultid="43069" />
                    <RANKING order="35" place="35" resultid="43128" />
                    <RANKING order="36" place="36" resultid="43013" />
                    <RANKING order="37" place="37" resultid="43816" />
                    <RANKING order="38" place="38" resultid="43488" />
                    <RANKING order="39" place="39" resultid="43324" />
                    <RANKING order="40" place="40" resultid="43880" />
                    <RANKING order="41" place="41" resultid="43350" />
                    <RANKING order="42" place="42" resultid="42493" />
                    <RANKING order="43" place="43" resultid="43810" />
                    <RANKING order="44" place="44" resultid="43483" />
                    <RANKING order="45" place="45" resultid="43451" />
                    <RANKING order="46" place="46" resultid="43182" />
                    <RANKING order="47" place="-1" resultid="41534" />
                    <RANKING order="48" place="-1" resultid="41828" />
                    <RANKING order="49" place="-1" resultid="42049" />
                    <RANKING order="50" place="-1" resultid="41652" />
                    <RANKING order="51" place="-1" resultid="41955" />
                    <RANKING order="52" place="-1" resultid="43984" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45079" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45080" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="45081" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="45082" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="45083" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="45084" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="45085" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2173" gender="F" number="3" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45156" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42330" />
                    <RANKING order="2" place="2" resultid="42356" />
                    <RANKING order="3" place="-1" resultid="43295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45157" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43079" />
                    <RANKING order="2" place="2" resultid="41541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45158" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45159" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43334" />
                    <RANKING order="2" place="2" resultid="43044" />
                    <RANKING order="3" place="-1" resultid="43526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45160" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43239" />
                    <RANKING order="2" place="2" resultid="43195" />
                    <RANKING order="3" place="3" resultid="42029" />
                    <RANKING order="4" place="4" resultid="43211" />
                    <RANKING order="5" place="5" resultid="41813" />
                    <RANKING order="6" place="-1" resultid="43180" />
                    <RANKING order="7" place="-1" resultid="43768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45161" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42044" />
                    <RANKING order="2" place="2" resultid="42241" />
                    <RANKING order="3" place="3" resultid="43900" />
                    <RANKING order="4" place="-1" resultid="41961" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45162" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42967" />
                    <RANKING order="2" place="2" resultid="43876" />
                    <RANKING order="3" place="3" resultid="42408" />
                    <RANKING order="4" place="-1" resultid="42070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45163" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43848" />
                    <RANKING order="2" place="2" resultid="43289" />
                    <RANKING order="3" place="3" resultid="43646" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45164" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="43954" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45165" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="43225" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45166" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45167" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45168" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45169" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45171" agemax="-1" agemin="-1" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43079" />
                    <RANKING order="2" place="2" resultid="42330" />
                    <RANKING order="3" place="3" resultid="42356" />
                    <RANKING order="4" place="4" resultid="42044" />
                    <RANKING order="5" place="5" resultid="41541" />
                    <RANKING order="6" place="6" resultid="43239" />
                    <RANKING order="7" place="7" resultid="42967" />
                    <RANKING order="8" place="8" resultid="43195" />
                    <RANKING order="9" place="9" resultid="43246" />
                    <RANKING order="10" place="10" resultid="43876" />
                    <RANKING order="11" place="11" resultid="43334" />
                    <RANKING order="12" place="12" resultid="43044" />
                    <RANKING order="13" place="13" resultid="42241" />
                    <RANKING order="14" place="14" resultid="43900" />
                    <RANKING order="15" place="15" resultid="42029" />
                    <RANKING order="16" place="16" resultid="43848" />
                    <RANKING order="17" place="17" resultid="42408" />
                    <RANKING order="18" place="18" resultid="43289" />
                    <RANKING order="19" place="19" resultid="43211" />
                    <RANKING order="20" place="20" resultid="43646" />
                    <RANKING order="21" place="21" resultid="41813" />
                    <RANKING order="22" place="-1" resultid="42070" />
                    <RANKING order="23" place="-1" resultid="43295" />
                    <RANKING order="24" place="-1" resultid="43180" />
                    <RANKING order="25" place="-1" resultid="43225" />
                    <RANKING order="26" place="-1" resultid="43526" />
                    <RANKING order="27" place="-1" resultid="43768" />
                    <RANKING order="28" place="-1" resultid="43954" />
                    <RANKING order="29" place="-1" resultid="41961" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45086" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45087" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="45088" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="45089" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2622" gender="M" number="4" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45187" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42683" />
                    <RANKING order="2" place="2" resultid="43083" />
                    <RANKING order="3" place="3" resultid="43484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45188" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43929" />
                    <RANKING order="2" place="2" resultid="42011" />
                    <RANKING order="3" place="3" resultid="43684" />
                    <RANKING order="4" place="4" resultid="42016" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45189" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43820" />
                    <RANKING order="2" place="2" resultid="42229" />
                    <RANKING order="3" place="3" resultid="43806" />
                    <RANKING order="4" place="4" resultid="42053" />
                    <RANKING order="5" place="5" resultid="43790" />
                    <RANKING order="6" place="6" resultid="41645" />
                    <RANKING order="7" place="7" resultid="43406" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45190" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42988" />
                    <RANKING order="2" place="2" resultid="44018" />
                    <RANKING order="3" place="3" resultid="42065" />
                    <RANKING order="4" place="4" resultid="43713" />
                    <RANKING order="5" place="-1" resultid="42188" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45191" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41807" />
                    <RANKING order="2" place="2" resultid="41737" />
                    <RANKING order="3" place="3" resultid="41864" />
                    <RANKING order="4" place="4" resultid="42828" />
                    <RANKING order="5" place="-1" resultid="43441" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45192" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42982" />
                    <RANKING order="2" place="2" resultid="42474" />
                    <RANKING order="3" place="3" resultid="43320" />
                    <RANKING order="4" place="4" resultid="42211" />
                    <RANKING order="5" place="5" resultid="42861" />
                    <RANKING order="6" place="6" resultid="41626" />
                    <RANKING order="7" place="7" resultid="43184" />
                    <RANKING order="8" place="8" resultid="43762" />
                    <RANKING order="9" place="9" resultid="43837" />
                    <RANKING order="10" place="-1" resultid="42855" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45193" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43204" />
                    <RANKING order="2" place="2" resultid="42223" />
                    <RANKING order="3" place="3" resultid="43014" />
                    <RANKING order="4" place="4" resultid="41892" />
                    <RANKING order="5" place="5" resultid="42144" />
                    <RANKING order="6" place="6" resultid="43962" />
                    <RANKING order="7" place="7" resultid="42437" />
                    <RANKING order="8" place="-1" resultid="41535" />
                    <RANKING order="9" place="-1" resultid="42978" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45194" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43213" />
                    <RANKING order="2" place="2" resultid="43489" />
                    <RANKING order="3" place="3" resultid="43452" />
                    <RANKING order="4" place="4" resultid="42126" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45195" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42099" />
                    <RANKING order="2" place="2" resultid="43263" />
                    <RANKING order="3" place="3" resultid="41699" />
                    <RANKING order="4" place="4" resultid="42150" />
                    <RANKING order="5" place="5" resultid="43493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45196" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42413" />
                    <RANKING order="2" place="2" resultid="41870" />
                    <RANKING order="3" place="3" resultid="43357" />
                    <RANKING order="4" place="4" resultid="41676" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45197" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41664" />
                    <RANKING order="2" place="2" resultid="43540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45198" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45199" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45200" agemax="94" agemin="90">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="41850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45201" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43929" />
                    <RANKING order="2" place="2" resultid="43820" />
                    <RANKING order="3" place="3" resultid="42011" />
                    <RANKING order="4" place="4" resultid="42229" />
                    <RANKING order="5" place="5" resultid="42988" />
                    <RANKING order="6" place="6" resultid="43684" />
                    <RANKING order="7" place="7" resultid="44018" />
                    <RANKING order="8" place="8" resultid="43204" />
                    <RANKING order="9" place="9" resultid="43806" />
                    <RANKING order="10" place="10" resultid="42982" />
                    <RANKING order="11" place="11" resultid="42683" />
                    <RANKING order="12" place="12" resultid="42223" />
                    <RANKING order="13" place="13" resultid="43083" />
                    <RANKING order="14" place="14" resultid="42474" />
                    <RANKING order="15" place="15" resultid="41807" />
                    <RANKING order="16" place="16" resultid="43213" />
                    <RANKING order="17" place="17" resultid="43320" />
                    <RANKING order="18" place="18" resultid="42053" />
                    <RANKING order="19" place="19" resultid="41737" />
                    <RANKING order="20" place="20" resultid="42065" />
                    <RANKING order="21" place="21" resultid="43713" />
                    <RANKING order="22" place="22" resultid="42016" />
                    <RANKING order="23" place="23" resultid="42211" />
                    <RANKING order="24" place="24" resultid="41864" />
                    <RANKING order="25" place="25" resultid="42828" />
                    <RANKING order="26" place="26" resultid="42861" />
                    <RANKING order="27" place="27" resultid="41626" />
                    <RANKING order="28" place="28" resultid="43184" />
                    <RANKING order="29" place="29" resultid="42099" />
                    <RANKING order="30" place="30" resultid="43790" />
                    <RANKING order="31" place="31" resultid="43762" />
                    <RANKING order="32" place="32" resultid="43837" />
                    <RANKING order="33" place="33" resultid="41645" />
                    <RANKING order="34" place="34" resultid="43263" />
                    <RANKING order="35" place="35" resultid="43014" />
                    <RANKING order="36" place="36" resultid="41892" />
                    <RANKING order="37" place="37" resultid="42144" />
                    <RANKING order="38" place="38" resultid="43484" />
                    <RANKING order="39" place="39" resultid="43406" />
                    <RANKING order="40" place="40" resultid="41664" />
                    <RANKING order="41" place="41" resultid="43962" />
                    <RANKING order="42" place="42" resultid="41699" />
                    <RANKING order="43" place="43" resultid="42413" />
                    <RANKING order="44" place="44" resultid="42437" />
                    <RANKING order="45" place="45" resultid="43489" />
                    <RANKING order="46" place="46" resultid="41870" />
                    <RANKING order="47" place="47" resultid="43452" />
                    <RANKING order="48" place="48" resultid="42150" />
                    <RANKING order="49" place="49" resultid="43357" />
                    <RANKING order="50" place="50" resultid="43540" />
                    <RANKING order="51" place="51" resultid="41676" />
                    <RANKING order="52" place="52" resultid="43493" />
                    <RANKING order="53" place="53" resultid="42126" />
                    <RANKING order="54" place="54" resultid="41904" />
                    <RANKING order="55" place="-1" resultid="42188" />
                    <RANKING order="56" place="-1" resultid="41535" />
                    <RANKING order="57" place="-1" resultid="41850" />
                    <RANKING order="58" place="-1" resultid="42855" />
                    <RANKING order="59" place="-1" resultid="42978" />
                    <RANKING order="60" place="-1" resultid="43441" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="44872" daytime="13:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="44873" daytime="13:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="44874" daytime="14:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="44875" daytime="14:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="44876" daytime="14:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="44877" daytime="14:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="44878" daytime="14:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="44879" daytime="14:25" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2203" gender="F" number="5" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45140" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42782" />
                    <RANKING order="2" place="2" resultid="42452" />
                    <RANKING order="3" place="3" resultid="42736" />
                    <RANKING order="4" place="4" resultid="42156" />
                    <RANKING order="5" place="5" resultid="43296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45141" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="45142" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41993" />
                    <RANKING order="2" place="2" resultid="42420" />
                    <RANKING order="3" place="3" resultid="43778" />
                    <RANKING order="4" place="4" resultid="42235" />
                    <RANKING order="5" place="5" resultid="43708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45143" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43843" />
                    <RANKING order="2" place="2" resultid="43904" />
                    <RANKING order="3" place="3" resultid="43045" />
                    <RANKING order="4" place="4" resultid="43335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45144" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41974" />
                    <RANKING order="2" place="2" resultid="43196" />
                    <RANKING order="3" place="3" resultid="42713" />
                    <RANKING order="4" place="4" resultid="43456" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45145" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43429" />
                    <RANKING order="2" place="2" resultid="41935" />
                    <RANKING order="3" place="-1" resultid="41710" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45146" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43435" />
                    <RANKING order="2" place="2" resultid="42132" />
                    <RANKING order="3" place="3" resultid="43328" />
                    <RANKING order="4" place="4" resultid="42205" />
                    <RANKING order="5" place="5" resultid="43235" />
                    <RANKING order="6" place="-1" resultid="42138" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45147" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42807" />
                    <RANKING order="2" place="2" resultid="41886" />
                    <RANKING order="3" place="-1" resultid="43570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45148" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45149" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="45150" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45151" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45152" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45153" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45154" agemax="94" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42782" />
                    <RANKING order="2" place="2" resultid="42452" />
                    <RANKING order="3" place="3" resultid="42736" />
                    <RANKING order="4" place="4" resultid="41993" />
                    <RANKING order="5" place="5" resultid="43843" />
                    <RANKING order="6" place="6" resultid="42156" />
                    <RANKING order="7" place="7" resultid="42420" />
                    <RANKING order="8" place="8" resultid="43435" />
                    <RANKING order="9" place="9" resultid="43778" />
                    <RANKING order="10" place="10" resultid="42132" />
                    <RANKING order="11" place="11" resultid="43904" />
                    <RANKING order="12" place="12" resultid="41974" />
                    <RANKING order="13" place="13" resultid="43328" />
                    <RANKING order="14" place="14" resultid="43429" />
                    <RANKING order="15" place="15" resultid="43296" />
                    <RANKING order="16" place="16" resultid="42235" />
                    <RANKING order="17" place="17" resultid="41935" />
                    <RANKING order="18" place="18" resultid="42205" />
                    <RANKING order="19" place="19" resultid="43196" />
                    <RANKING order="20" place="20" resultid="42713" />
                    <RANKING order="21" place="21" resultid="43708" />
                    <RANKING order="22" place="22" resultid="43045" />
                    <RANKING order="23" place="23" resultid="43335" />
                    <RANKING order="24" place="24" resultid="43235" />
                    <RANKING order="25" place="25" resultid="43456" />
                    <RANKING order="26" place="26" resultid="41881" />
                    <RANKING order="27" place="27" resultid="42807" />
                    <RANKING order="28" place="28" resultid="41886" />
                    <RANKING order="29" place="-1" resultid="41710" />
                    <RANKING order="30" place="-1" resultid="42138" />
                    <RANKING order="31" place="-1" resultid="43570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45155" agemax="-1" agemin="-1" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42782" />
                    <RANKING order="2" place="2" resultid="42452" />
                    <RANKING order="3" place="3" resultid="42736" />
                    <RANKING order="4" place="4" resultid="41993" />
                    <RANKING order="5" place="5" resultid="43843" />
                    <RANKING order="6" place="6" resultid="42156" />
                    <RANKING order="7" place="7" resultid="42420" />
                    <RANKING order="8" place="8" resultid="43435" />
                    <RANKING order="9" place="9" resultid="43778" />
                    <RANKING order="10" place="10" resultid="42132" />
                    <RANKING order="11" place="11" resultid="43904" />
                    <RANKING order="12" place="12" resultid="41974" />
                    <RANKING order="13" place="13" resultid="43328" />
                    <RANKING order="14" place="14" resultid="43429" />
                    <RANKING order="15" place="15" resultid="43296" />
                    <RANKING order="16" place="16" resultid="42235" />
                    <RANKING order="17" place="17" resultid="41935" />
                    <RANKING order="18" place="18" resultid="42205" />
                    <RANKING order="19" place="19" resultid="43196" />
                    <RANKING order="20" place="20" resultid="42713" />
                    <RANKING order="21" place="21" resultid="43708" />
                    <RANKING order="22" place="22" resultid="43045" />
                    <RANKING order="23" place="23" resultid="43335" />
                    <RANKING order="24" place="24" resultid="43235" />
                    <RANKING order="25" place="25" resultid="43456" />
                    <RANKING order="26" place="26" resultid="41881" />
                    <RANKING order="27" place="27" resultid="42807" />
                    <RANKING order="28" place="28" resultid="41886" />
                    <RANKING order="29" place="-1" resultid="41710" />
                    <RANKING order="30" place="-1" resultid="42138" />
                    <RANKING order="31" place="-1" resultid="43570" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="44880" daytime="14:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="44881" daytime="14:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="44882" daytime="14:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="44883" daytime="14:40" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2537" gender="M" number="6" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45172" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42700" />
                    <RANKING order="2" place="2" resultid="43339" />
                    <RANKING order="3" place="3" resultid="42674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45173" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42017" />
                    <RANKING order="2" place="-1" resultid="42022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45174" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42058" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45175" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43942" />
                    <RANKING order="2" place="2" resultid="41908" />
                    <RANKING order="3" place="3" resultid="41836" />
                    <RANKING order="4" place="-1" resultid="42246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45176" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41842" />
                    <RANKING order="2" place="2" resultid="42194" />
                    <RANKING order="3" place="3" resultid="43377" />
                    <RANKING order="4" place="4" resultid="41865" />
                    <RANKING order="5" place="5" resultid="43418" />
                    <RANKING order="6" place="6" resultid="43325" />
                    <RANKING order="7" place="-1" resultid="43994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45177" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43314" />
                    <RANKING order="2" place="2" resultid="42217" />
                    <RANKING order="3" place="3" resultid="43321" />
                    <RANKING order="4" place="4" resultid="42719" />
                    <RANKING order="5" place="5" resultid="43502" />
                    <RANKING order="6" place="6" resultid="43831" />
                    <RANKING order="7" place="7" resultid="43049" />
                    <RANKING order="8" place="-1" resultid="42109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45178" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42224" />
                    <RANKING order="2" place="2" resultid="43800" />
                    <RANKING order="3" place="3" resultid="43057" />
                    <RANKING order="4" place="4" resultid="41893" />
                    <RANKING order="5" place="5" resultid="41858" />
                    <RANKING order="6" place="6" resultid="43963" />
                    <RANKING order="7" place="-1" resultid="43923" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45179" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42037" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45180" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43264" />
                    <RANKING order="2" place="2" resultid="43129" />
                    <RANKING order="3" place="3" resultid="43025" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45181" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="45182" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43580" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45183" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45184" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45185" agemax="94" agemin="90">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="41851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45186" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42700" />
                    <RANKING order="2" place="2" resultid="41842" />
                    <RANKING order="3" place="3" resultid="43314" />
                    <RANKING order="4" place="4" resultid="42194" />
                    <RANKING order="5" place="5" resultid="42217" />
                    <RANKING order="6" place="6" resultid="43339" />
                    <RANKING order="7" place="7" resultid="43942" />
                    <RANKING order="8" place="8" resultid="42674" />
                    <RANKING order="9" place="9" resultid="43321" />
                    <RANKING order="10" place="10" resultid="42224" />
                    <RANKING order="11" place="11" resultid="43800" />
                    <RANKING order="12" place="12" resultid="41908" />
                    <RANKING order="13" place="13" resultid="41836" />
                    <RANKING order="14" place="14" resultid="43377" />
                    <RANKING order="15" place="15" resultid="42058" />
                    <RANKING order="16" place="16" resultid="42017" />
                    <RANKING order="17" place="17" resultid="42719" />
                    <RANKING order="18" place="18" resultid="41865" />
                    <RANKING order="19" place="19" resultid="43057" />
                    <RANKING order="20" place="20" resultid="41893" />
                    <RANKING order="21" place="21" resultid="43502" />
                    <RANKING order="22" place="22" resultid="41858" />
                    <RANKING order="23" place="23" resultid="43418" />
                    <RANKING order="24" place="24" resultid="43831" />
                    <RANKING order="25" place="25" resultid="43264" />
                    <RANKING order="26" place="26" resultid="43129" />
                    <RANKING order="27" place="27" resultid="42037" />
                    <RANKING order="28" place="28" resultid="43049" />
                    <RANKING order="29" place="29" resultid="43025" />
                    <RANKING order="30" place="30" resultid="43963" />
                    <RANKING order="31" place="31" resultid="43325" />
                    <RANKING order="32" place="32" resultid="43580" />
                    <RANKING order="33" place="-1" resultid="41851" />
                    <RANKING order="34" place="-1" resultid="42022" />
                    <RANKING order="35" place="-1" resultid="42109" />
                    <RANKING order="36" place="-1" resultid="42246" />
                    <RANKING order="37" place="-1" resultid="43923" />
                    <RANKING order="38" place="-1" resultid="43994" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="44884" daytime="14:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="44885" daytime="14:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="44886" daytime="14:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="44887" daytime="14:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="44888" daytime="15:00" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2021-07-09" daytime="15:30" endtime="19:37" name="1ª Jornada-2ª sessão" number="2" warmupfrom="08:00" warmupuntil="09:15">
          <EVENTS>
            <EVENT eventid="2338" daytime="15:30" gender="F" number="7" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45267" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42499" />
                    <RANKING order="2" place="2" resultid="42783" />
                    <RANKING order="3" place="3" resultid="42737" />
                    <RANKING order="4" place="4" resultid="44028" />
                    <RANKING order="5" place="5" resultid="43008" />
                    <RANKING order="6" place="6" resultid="44033" />
                    <RANKING order="7" place="7" resultid="43297" />
                    <RANKING order="8" place="-1" resultid="42350" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45268" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41723" />
                    <RANKING order="2" place="2" resultid="43661" />
                    <RANKING order="3" place="3" resultid="42076" />
                    <RANKING order="4" place="-1" resultid="42200" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45269" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="41769" />
                    <RANKING order="2" place="-1" resultid="41523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45270" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43844" />
                    <RANKING order="2" place="2" resultid="43037" />
                    <RANKING order="3" place="3" resultid="42731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45271" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43277" />
                    <RANKING order="2" place="2" resultid="41971" />
                    <RANKING order="3" place="3" resultid="41814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45272" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43300" />
                    <RANKING order="2" place="2" resultid="42174" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45273" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42133" />
                    <RANKING order="2" place="2" resultid="41854" />
                    <RANKING order="3" place="3" resultid="42206" />
                    <RANKING order="4" place="4" resultid="43756" />
                    <RANKING order="5" place="5" resultid="43123" />
                    <RANKING order="6" place="6" resultid="41756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45274" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43849" />
                    <RANKING order="2" place="2" resultid="41744" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45275" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="45276" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="45277" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45278" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45279" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45280" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45281" agemax="-1" agemin="-1" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42499" />
                    <RANKING order="2" place="2" resultid="42783" />
                    <RANKING order="3" place="3" resultid="41723" />
                    <RANKING order="4" place="4" resultid="43661" />
                    <RANKING order="5" place="5" resultid="43844" />
                    <RANKING order="6" place="6" resultid="43277" />
                    <RANKING order="7" place="7" resultid="42737" />
                    <RANKING order="8" place="8" resultid="43037" />
                    <RANKING order="9" place="9" resultid="42076" />
                    <RANKING order="10" place="10" resultid="44028" />
                    <RANKING order="11" place="11" resultid="43300" />
                    <RANKING order="12" place="12" resultid="43008" />
                    <RANKING order="13" place="13" resultid="42133" />
                    <RANKING order="14" place="14" resultid="42731" />
                    <RANKING order="15" place="15" resultid="41971" />
                    <RANKING order="16" place="16" resultid="44033" />
                    <RANKING order="17" place="17" resultid="41854" />
                    <RANKING order="18" place="18" resultid="43297" />
                    <RANKING order="19" place="19" resultid="42206" />
                    <RANKING order="20" place="20" resultid="42174" />
                    <RANKING order="21" place="21" resultid="43849" />
                    <RANKING order="22" place="22" resultid="43756" />
                    <RANKING order="23" place="23" resultid="43123" />
                    <RANKING order="24" place="24" resultid="41744" />
                    <RANKING order="25" place="25" resultid="41756" />
                    <RANKING order="26" place="26" resultid="41814" />
                    <RANKING order="27" place="-1" resultid="41769" />
                    <RANKING order="28" place="-1" resultid="42200" />
                    <RANKING order="29" place="-1" resultid="42350" />
                    <RANKING order="30" place="-1" resultid="41523" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="44889" daytime="15:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="44890" daytime="15:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="44891" daytime="15:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="44892" daytime="15:35" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2682" daytime="15:40" gender="M" number="8" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45237" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42323" />
                    <RANKING order="2" place="2" resultid="42818" />
                    <RANKING order="3" place="3" resultid="42701" />
                    <RANKING order="4" place="4" resultid="43933" />
                    <RANKING order="5" place="5" resultid="42834" />
                    <RANKING order="6" place="6" resultid="42795" />
                    <RANKING order="7" place="7" resultid="42374" />
                    <RANKING order="8" place="8" resultid="42865" />
                    <RANKING order="9" place="9" resultid="41732" />
                    <RANKING order="10" place="10" resultid="42675" />
                    <RANKING order="11" place="11" resultid="43703" />
                    <RANKING order="12" place="12" resultid="42684" />
                    <RANKING order="13" place="-1" resultid="42338" />
                    <RANKING order="14" place="-1" resultid="43001" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45238" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43741" />
                    <RANKING order="2" place="2" resultid="43818" />
                    <RANKING order="3" place="3" resultid="42709" />
                    <RANKING order="4" place="4" resultid="43783" />
                    <RANKING order="5" place="5" resultid="41949" />
                    <RANKING order="6" place="-1" resultid="41529" />
                    <RANKING order="7" place="-1" resultid="43858" />
                    <RANKING order="8" place="-1" resultid="43952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45239" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42771" />
                    <RANKING order="2" place="2" resultid="43917" />
                    <RANKING order="3" place="3" resultid="42483" />
                    <RANKING order="4" place="4" resultid="42230" />
                    <RANKING order="5" place="5" resultid="43699" />
                    <RANKING order="6" place="6" resultid="41646" />
                    <RANKING order="7" place="7" resultid="43791" />
                    <RANKING order="8" place="8" resultid="43718" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45240" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43363" />
                    <RANKING order="2" place="2" resultid="42763" />
                    <RANKING order="3" place="3" resultid="44019" />
                    <RANKING order="4" place="4" resultid="42189" />
                    <RANKING order="5" place="5" resultid="43694" />
                    <RANKING order="6" place="-1" resultid="44001" />
                    <RANKING order="7" place="-1" resultid="41518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45241" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43586" />
                    <RANKING order="2" place="2" resultid="42195" />
                    <RANKING order="3" place="3" resultid="41843" />
                    <RANKING order="4" place="4" resultid="41790" />
                    <RANKING order="5" place="5" resultid="42961" />
                    <RANKING order="6" place="6" resultid="43546" />
                    <RANKING order="7" place="7" resultid="41808" />
                    <RANKING order="8" place="8" resultid="42171" />
                    <RANKING order="9" place="9" resultid="42832" />
                    <RANKING order="10" place="10" resultid="43989" />
                    <RANKING order="11" place="11" resultid="43445" />
                    <RANKING order="12" place="-1" resultid="43854" />
                    <RANKING order="13" place="-1" resultid="43985" />
                    <RANKING order="14" place="-1" resultid="43995" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45242" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43389" />
                    <RANKING order="2" place="2" resultid="41632" />
                    <RANKING order="3" place="3" resultid="43315" />
                    <RANKING order="4" place="4" resultid="43259" />
                    <RANKING order="5" place="5" resultid="43382" />
                    <RANKING order="6" place="6" resultid="42212" />
                    <RANKING order="7" place="7" resultid="42720" />
                    <RANKING order="8" place="8" resultid="44024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45243" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43563" />
                    <RANKING order="2" place="2" resultid="43801" />
                    <RANKING order="3" place="3" resultid="43070" />
                    <RANKING order="4" place="-1" resultid="43619" />
                    <RANKING order="5" place="-1" resultid="43508" />
                    <RANKING order="6" place="-1" resultid="43924" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45244" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43513" />
                    <RANKING order="2" place="2" resultid="43214" />
                    <RANKING order="3" place="3" resultid="42115" />
                    <RANKING order="4" place="4" resultid="43881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45245" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43019" />
                    <RANKING order="2" place="2" resultid="43494" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45246" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41659" />
                    <RANKING order="2" place="2" resultid="42743" />
                    <RANKING order="3" place="3" resultid="43358" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45247" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45248" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45249" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45250" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45251" agemax="94" agemin="25" name="Absolutos">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43741" />
                    <RANKING order="2" place="2" resultid="42323" />
                    <RANKING order="3" place="3" resultid="42818" />
                    <RANKING order="4" place="4" resultid="43818" />
                    <RANKING order="5" place="5" resultid="42701" />
                    <RANKING order="6" place="6" resultid="42771" />
                    <RANKING order="7" place="7" resultid="43933" />
                    <RANKING order="8" place="8" resultid="42834" />
                    <RANKING order="9" place="9" resultid="43917" />
                    <RANKING order="10" place="10" resultid="42483" />
                    <RANKING order="11" place="11" resultid="43586" />
                    <RANKING order="12" place="12" resultid="42230" />
                    <RANKING order="13" place="13" resultid="43389" />
                    <RANKING order="14" place="14" resultid="42195" />
                    <RANKING order="15" place="15" resultid="42795" />
                    <RANKING order="16" place="16" resultid="41632" />
                    <RANKING order="17" place="17" resultid="42374" />
                    <RANKING order="18" place="18" resultid="41843" />
                    <RANKING order="19" place="18" resultid="42709" />
                    <RANKING order="20" place="18" resultid="43363" />
                    <RANKING order="21" place="21" resultid="42865" />
                    <RANKING order="22" place="22" resultid="43315" />
                    <RANKING order="23" place="23" resultid="41732" />
                    <RANKING order="24" place="24" resultid="41790" />
                    <RANKING order="25" place="25" resultid="43259" />
                    <RANKING order="26" place="26" resultid="43563" />
                    <RANKING order="27" place="27" resultid="42961" />
                    <RANKING order="28" place="28" resultid="42763" />
                    <RANKING order="29" place="29" resultid="42675" />
                    <RANKING order="30" place="30" resultid="43699" />
                    <RANKING order="31" place="31" resultid="43382" />
                    <RANKING order="32" place="32" resultid="44019" />
                    <RANKING order="33" place="33" resultid="42189" />
                    <RANKING order="34" place="34" resultid="43783" />
                    <RANKING order="35" place="35" resultid="41949" />
                    <RANKING order="36" place="36" resultid="43546" />
                    <RANKING order="37" place="37" resultid="41808" />
                    <RANKING order="38" place="38" resultid="43513" />
                    <RANKING order="39" place="39" resultid="43703" />
                    <RANKING order="40" place="40" resultid="42684" />
                    <RANKING order="41" place="41" resultid="43801" />
                    <RANKING order="42" place="42" resultid="42212" />
                    <RANKING order="43" place="43" resultid="43214" />
                    <RANKING order="44" place="44" resultid="42115" />
                    <RANKING order="45" place="45" resultid="42171" />
                    <RANKING order="46" place="46" resultid="42832" />
                    <RANKING order="47" place="47" resultid="42720" />
                    <RANKING order="48" place="48" resultid="44024" />
                    <RANKING order="49" place="49" resultid="43989" />
                    <RANKING order="50" place="50" resultid="41646" />
                    <RANKING order="51" place="51" resultid="43791" />
                    <RANKING order="52" place="52" resultid="43718" />
                    <RANKING order="53" place="53" resultid="43445" />
                    <RANKING order="54" place="54" resultid="43070" />
                    <RANKING order="55" place="55" resultid="41659" />
                    <RANKING order="56" place="56" resultid="43694" />
                    <RANKING order="57" place="57" resultid="43019" />
                    <RANKING order="58" place="58" resultid="42743" />
                    <RANKING order="59" place="59" resultid="43881" />
                    <RANKING order="60" place="60" resultid="43358" />
                    <RANKING order="61" place="61" resultid="43494" />
                    <RANKING order="62" place="-1" resultid="43619" />
                    <RANKING order="63" place="-1" resultid="41529" />
                    <RANKING order="64" place="-1" resultid="42338" />
                    <RANKING order="65" place="-1" resultid="43001" />
                    <RANKING order="66" place="-1" resultid="43508" />
                    <RANKING order="67" place="-1" resultid="43854" />
                    <RANKING order="68" place="-1" resultid="43858" />
                    <RANKING order="69" place="-1" resultid="43924" />
                    <RANKING order="70" place="-1" resultid="43952" />
                    <RANKING order="71" place="-1" resultid="44001" />
                    <RANKING order="72" place="-1" resultid="41518" />
                    <RANKING order="73" place="-1" resultid="43985" />
                    <RANKING order="74" place="-1" resultid="43995" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="44893" daytime="15:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="44894" daytime="15:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="44895" daytime="15:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="44896" daytime="15:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="44897" daytime="15:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="44898" daytime="15:50" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="44899" daytime="15:50" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="44900" daytime="15:55" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="44901" daytime="15:55" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2278" daytime="15:55" gender="F" number="9" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45282" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43667" />
                    <RANKING order="2" place="2" resultid="42500" />
                    <RANKING order="3" place="3" resultid="42453" />
                    <RANKING order="4" place="4" resultid="42351" />
                    <RANKING order="5" place="5" resultid="42463" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45283" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42077" />
                    <RANKING order="2" place="2" resultid="41542" />
                    <RANKING order="3" place="-1" resultid="42201" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45284" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="41524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45285" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43527" />
                    <RANKING order="2" place="2" resultid="42696" />
                    <RANKING order="3" place="3" resultid="43905" />
                    <RANKING order="4" place="4" resultid="43038" />
                    <RANKING order="5" place="5" resultid="43398" />
                    <RANKING order="6" place="6" resultid="41546" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45286" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42082" />
                    <RANKING order="2" place="2" resultid="43278" />
                    <RANKING order="3" place="3" resultid="42714" />
                    <RANKING order="4" place="4" resultid="42839" />
                    <RANKING order="5" place="-1" resultid="41940" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45287" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43221" />
                    <RANKING order="2" place="2" resultid="43430" />
                    <RANKING order="3" place="3" resultid="43679" />
                    <RANKING order="4" place="-1" resultid="41711" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45288" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42139" />
                    <RANKING order="2" place="2" resultid="43436" />
                    <RANKING order="3" place="3" resultid="41919" />
                    <RANKING order="4" place="4" resultid="43329" />
                    <RANKING order="5" place="5" resultid="43124" />
                    <RANKING order="6" place="6" resultid="42690" />
                    <RANKING order="7" place="7" resultid="43650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45289" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="43571" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45290" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45291" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="45292" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45293" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45294" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45295" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45296" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43667" />
                    <RANKING order="2" place="2" resultid="42500" />
                    <RANKING order="3" place="3" resultid="42453" />
                    <RANKING order="4" place="4" resultid="42082" />
                    <RANKING order="5" place="5" resultid="43278" />
                    <RANKING order="6" place="6" resultid="43221" />
                    <RANKING order="7" place="7" resultid="42351" />
                    <RANKING order="8" place="8" resultid="43527" />
                    <RANKING order="9" place="9" resultid="42696" />
                    <RANKING order="10" place="10" resultid="42139" />
                    <RANKING order="11" place="11" resultid="43905" />
                    <RANKING order="12" place="12" resultid="43038" />
                    <RANKING order="13" place="13" resultid="42077" />
                    <RANKING order="14" place="14" resultid="42463" />
                    <RANKING order="15" place="15" resultid="43436" />
                    <RANKING order="16" place="16" resultid="43398" />
                    <RANKING order="17" place="17" resultid="41542" />
                    <RANKING order="18" place="18" resultid="41919" />
                    <RANKING order="19" place="19" resultid="43329" />
                    <RANKING order="20" place="20" resultid="43430" />
                    <RANKING order="21" place="21" resultid="43124" />
                    <RANKING order="22" place="22" resultid="41546" />
                    <RANKING order="23" place="23" resultid="43679" />
                    <RANKING order="24" place="24" resultid="42714" />
                    <RANKING order="25" place="25" resultid="42690" />
                    <RANKING order="26" place="26" resultid="42839" />
                    <RANKING order="27" place="27" resultid="43650" />
                    <RANKING order="28" place="28" resultid="43534" />
                    <RANKING order="29" place="-1" resultid="41711" />
                    <RANKING order="30" place="-1" resultid="42201" />
                    <RANKING order="31" place="-1" resultid="43571" />
                    <RANKING order="32" place="-1" resultid="41524" />
                    <RANKING order="33" place="-1" resultid="41940" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="44902" daytime="15:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="44903" daytime="16:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="44904" daytime="16:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="44905" daytime="16:10" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2507" daytime="16:15" gender="M" number="10" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45252" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42324" />
                    <RANKING order="2" place="2" resultid="42813" />
                    <RANKING order="3" place="3" resultid="42369" />
                    <RANKING order="4" place="4" resultid="43485" />
                    <RANKING order="5" place="-1" resultid="42339" />
                    <RANKING order="6" place="-1" resultid="43737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45253" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43742" />
                    <RANKING order="2" place="2" resultid="42431" />
                    <RANKING order="3" place="3" resultid="43310" />
                    <RANKING order="4" place="4" resultid="43673" />
                    <RANKING order="5" place="5" resultid="43631" />
                    <RANKING order="6" place="-1" resultid="42023" />
                    <RANKING order="7" place="-1" resultid="43859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45254" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43075" />
                    <RANKING order="2" place="2" resultid="42059" />
                    <RANKING order="3" place="3" resultid="43407" />
                    <RANKING order="4" place="-1" resultid="41829" />
                    <RANKING order="5" place="-1" resultid="43472" />
                    <RANKING order="6" place="-1" resultid="42468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45255" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42087" />
                    <RANKING order="2" place="2" resultid="43695" />
                    <RANKING order="3" place="-1" resultid="41519" />
                    <RANKING order="4" place="-1" resultid="41956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45256" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43174" />
                    <RANKING order="2" place="2" resultid="42196" />
                    <RANKING order="3" place="3" resultid="41966" />
                    <RANKING order="4" place="4" resultid="43547" />
                    <RANKING order="5" place="5" resultid="42094" />
                    <RANKING order="6" place="6" resultid="43690" />
                    <RANKING order="7" place="7" resultid="42959" />
                    <RANKING order="8" place="8" resultid="42829" />
                    <RANKING order="9" place="9" resultid="43446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45257" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41633" />
                    <RANKING order="2" place="2" resultid="43316" />
                    <RANKING order="3" place="3" resultid="43322" />
                    <RANKING order="4" place="4" resultid="42180" />
                    <RANKING order="5" place="5" resultid="42983" />
                    <RANKING order="6" place="6" resultid="43503" />
                    <RANKING order="7" place="7" resultid="43832" />
                    <RANKING order="8" place="8" resultid="43050" />
                    <RANKING order="9" place="-1" resultid="42110" />
                    <RANKING order="10" place="-1" resultid="42856" />
                    <RANKING order="11" place="-1" resultid="43590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45258" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43611" />
                    <RANKING order="2" place="2" resultid="41716" />
                    <RANKING order="3" place="3" resultid="43205" />
                    <RANKING order="4" place="4" resultid="43190" />
                    <RANKING order="5" place="-1" resultid="41536" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45259" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41685" />
                    <RANKING order="2" place="2" resultid="43520" />
                    <RANKING order="3" place="3" resultid="43490" />
                    <RANKING order="4" place="4" resultid="42038" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45260" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43130" />
                    <RANKING order="2" place="2" resultid="42749" />
                    <RANKING order="3" place="3" resultid="41762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45261" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41660" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45262" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41653" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45263" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45264" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45265" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45266" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43742" />
                    <RANKING order="2" place="2" resultid="42324" />
                    <RANKING order="3" place="3" resultid="42087" />
                    <RANKING order="4" place="4" resultid="43611" />
                    <RANKING order="5" place="5" resultid="43174" />
                    <RANKING order="6" place="6" resultid="42813" />
                    <RANKING order="7" place="7" resultid="41633" />
                    <RANKING order="8" place="8" resultid="42369" />
                    <RANKING order="9" place="9" resultid="42196" />
                    <RANKING order="10" place="10" resultid="43316" />
                    <RANKING order="11" place="11" resultid="42431" />
                    <RANKING order="12" place="12" resultid="43322" />
                    <RANKING order="13" place="13" resultid="43310" />
                    <RANKING order="14" place="14" resultid="41685" />
                    <RANKING order="15" place="15" resultid="43673" />
                    <RANKING order="16" place="16" resultid="41716" />
                    <RANKING order="17" place="17" resultid="41966" />
                    <RANKING order="18" place="18" resultid="43631" />
                    <RANKING order="19" place="19" resultid="43205" />
                    <RANKING order="20" place="20" resultid="43547" />
                    <RANKING order="21" place="21" resultid="42180" />
                    <RANKING order="22" place="22" resultid="42094" />
                    <RANKING order="23" place="23" resultid="43690" />
                    <RANKING order="24" place="24" resultid="42959" />
                    <RANKING order="25" place="25" resultid="43520" />
                    <RANKING order="26" place="26" resultid="43075" />
                    <RANKING order="27" place="27" resultid="42983" />
                    <RANKING order="28" place="28" resultid="41660" />
                    <RANKING order="29" place="29" resultid="42059" />
                    <RANKING order="30" place="30" resultid="43190" />
                    <RANKING order="31" place="31" resultid="42829" />
                    <RANKING order="32" place="32" resultid="43503" />
                    <RANKING order="33" place="33" resultid="43695" />
                    <RANKING order="34" place="34" resultid="43130" />
                    <RANKING order="35" place="35" resultid="42749" />
                    <RANKING order="36" place="36" resultid="43446" />
                    <RANKING order="37" place="37" resultid="43832" />
                    <RANKING order="38" place="38" resultid="43490" />
                    <RANKING order="39" place="39" resultid="43050" />
                    <RANKING order="40" place="40" resultid="41762" />
                    <RANKING order="41" place="41" resultid="43407" />
                    <RANKING order="42" place="42" resultid="42038" />
                    <RANKING order="43" place="43" resultid="41653" />
                    <RANKING order="44" place="44" resultid="43485" />
                    <RANKING order="45" place="-1" resultid="41536" />
                    <RANKING order="46" place="-1" resultid="41829" />
                    <RANKING order="47" place="-1" resultid="42023" />
                    <RANKING order="48" place="-1" resultid="42110" />
                    <RANKING order="49" place="-1" resultid="42856" />
                    <RANKING order="50" place="-1" resultid="43472" />
                    <RANKING order="51" place="-1" resultid="43590" />
                    <RANKING order="52" place="-1" resultid="43859" />
                    <RANKING order="53" place="-1" resultid="41519" />
                    <RANKING order="54" place="-1" resultid="41956" />
                    <RANKING order="55" place="-1" resultid="42339" />
                    <RANKING order="56" place="-1" resultid="42468" />
                    <RANKING order="57" place="-1" resultid="43737" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45090" daytime="16:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45091" daytime="16:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="45092" daytime="16:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="45093" daytime="16:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="45094" daytime="16:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="45095" daytime="16:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="45096" daytime="16:45" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2021-07-10" daytime="09:30" endtime="18:10" name="2ª Jornada-1ª sessão" number="3" warmupfrom="08:00" warmupuntil="09:15">
          <EVENTS>
            <EVENT eventid="2308" daytime="09:30" gender="F" number="11" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45614" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42784" />
                    <RANKING order="2" place="2" resultid="42157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45615" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45616" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42236" />
                    <RANKING order="2" place="2" resultid="43709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45617" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43845" />
                    <RANKING order="2" place="2" resultid="43399" />
                    <RANKING order="3" place="3" resultid="43336" />
                    <RANKING order="4" place="4" resultid="43046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45618" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42120" />
                    <RANKING order="2" place="2" resultid="43197" />
                    <RANKING order="3" place="3" resultid="42030" />
                    <RANKING order="4" place="4" resultid="43457" />
                    <RANKING order="5" place="-1" resultid="43828" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45619" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42045" />
                    <RANKING order="2" place="2" resultid="42458" />
                    <RANKING order="3" place="3" resultid="41936" />
                    <RANKING order="4" place="4" resultid="43054" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45620" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43437" />
                    <RANKING order="2" place="2" resultid="42134" />
                    <RANKING order="3" place="3" resultid="43330" />
                    <RANKING order="4" place="4" resultid="42207" />
                    <RANKING order="5" place="5" resultid="43236" />
                    <RANKING order="6" place="6" resultid="43477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45621" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="45622" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="45623" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="45624" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45625" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45626" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45627" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45628" agemax="-1" agemin="-1" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42784" />
                    <RANKING order="2" place="2" resultid="42120" />
                    <RANKING order="3" place="3" resultid="43845" />
                    <RANKING order="4" place="4" resultid="42442" />
                    <RANKING order="5" place="5" resultid="42157" />
                    <RANKING order="6" place="6" resultid="42045" />
                    <RANKING order="7" place="7" resultid="43437" />
                    <RANKING order="8" place="8" resultid="42458" />
                    <RANKING order="9" place="9" resultid="42134" />
                    <RANKING order="10" place="10" resultid="43330" />
                    <RANKING order="11" place="11" resultid="42236" />
                    <RANKING order="12" place="12" resultid="41936" />
                    <RANKING order="13" place="13" resultid="42207" />
                    <RANKING order="14" place="14" resultid="43197" />
                    <RANKING order="15" place="15" resultid="43399" />
                    <RANKING order="16" place="16" resultid="43336" />
                    <RANKING order="17" place="17" resultid="43709" />
                    <RANKING order="18" place="18" resultid="42030" />
                    <RANKING order="19" place="19" resultid="43046" />
                    <RANKING order="20" place="20" resultid="43236" />
                    <RANKING order="21" place="21" resultid="43457" />
                    <RANKING order="22" place="22" resultid="43054" />
                    <RANKING order="23" place="23" resultid="43477" />
                    <RANKING order="24" place="-1" resultid="43828" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="44913" daytime="09:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="44914" daytime="09:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="44915" daytime="09:45" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2218" daytime="09:50" gender="M" number="12" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45449" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43340" />
                    <RANKING order="2" place="-1" resultid="42788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45450" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42018" />
                    <RANKING order="2" place="-1" resultid="42024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45451" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43821" />
                    <RANKING order="2" place="2" resultid="43945" />
                    <RANKING order="3" place="3" resultid="42005" />
                    <RANKING order="4" place="4" resultid="42060" />
                    <RANKING order="5" place="5" resultid="43792" />
                    <RANKING order="6" place="6" resultid="43408" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45452" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43460" />
                    <RANKING order="2" place="2" resultid="41909" />
                    <RANKING order="3" place="-1" resultid="41750" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45453" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41844" />
                    <RANKING order="2" place="2" resultid="42197" />
                    <RANKING order="3" place="3" resultid="43531" />
                    <RANKING order="4" place="4" resultid="43419" />
                    <RANKING order="5" place="5" resultid="41866" />
                    <RANKING order="6" place="6" resultid="43447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45454" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42218" />
                    <RANKING order="2" place="2" resultid="42488" />
                    <RANKING order="3" place="3" resultid="41898" />
                    <RANKING order="4" place="4" resultid="43886" />
                    <RANKING order="5" place="5" resultid="43504" />
                    <RANKING order="6" place="6" resultid="42721" />
                    <RANKING order="7" place="-1" resultid="43833" />
                    <RANKING order="8" place="-1" resultid="42111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45455" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43345" />
                    <RANKING order="2" place="2" resultid="42225" />
                    <RANKING order="3" place="3" resultid="43802" />
                    <RANKING order="4" place="4" resultid="41859" />
                    <RANKING order="5" place="5" resultid="41999" />
                    <RANKING order="6" place="6" resultid="43015" />
                    <RANKING order="7" place="7" resultid="41670" />
                    <RANKING order="8" place="-1" resultid="43058" />
                    <RANKING order="9" place="-1" resultid="42165" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45456" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42973" />
                    <RANKING order="2" place="2" resultid="43882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45457" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41693" />
                    <RANKING order="2" place="2" resultid="43026" />
                    <RANKING order="3" place="3" resultid="42151" />
                    <RANKING order="4" place="-1" resultid="42100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45458" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="45459" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45460" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45461" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45462" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45463" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43821" />
                    <RANKING order="2" place="2" resultid="43945" />
                    <RANKING order="3" place="3" resultid="41844" />
                    <RANKING order="4" place="4" resultid="42973" />
                    <RANKING order="5" place="5" resultid="42005" />
                    <RANKING order="6" place="6" resultid="42197" />
                    <RANKING order="7" place="7" resultid="43340" />
                    <RANKING order="8" place="8" resultid="42218" />
                    <RANKING order="9" place="9" resultid="43345" />
                    <RANKING order="10" place="10" resultid="43460" />
                    <RANKING order="11" place="11" resultid="42488" />
                    <RANKING order="12" place="12" resultid="42225" />
                    <RANKING order="13" place="13" resultid="41909" />
                    <RANKING order="14" place="14" resultid="41693" />
                    <RANKING order="15" place="15" resultid="43802" />
                    <RANKING order="16" place="16" resultid="41898" />
                    <RANKING order="17" place="17" resultid="43886" />
                    <RANKING order="18" place="18" resultid="42060" />
                    <RANKING order="19" place="19" resultid="42018" />
                    <RANKING order="20" place="20" resultid="43504" />
                    <RANKING order="21" place="21" resultid="42721" />
                    <RANKING order="22" place="22" resultid="43531" />
                    <RANKING order="23" place="23" resultid="43419" />
                    <RANKING order="24" place="24" resultid="41859" />
                    <RANKING order="25" place="25" resultid="41866" />
                    <RANKING order="26" place="26" resultid="43792" />
                    <RANKING order="27" place="27" resultid="41999" />
                    <RANKING order="28" place="28" resultid="43015" />
                    <RANKING order="29" place="29" resultid="43408" />
                    <RANKING order="30" place="30" resultid="43882" />
                    <RANKING order="31" place="31" resultid="43447" />
                    <RANKING order="32" place="32" resultid="43026" />
                    <RANKING order="33" place="33" resultid="41670" />
                    <RANKING order="34" place="34" resultid="43581" />
                    <RANKING order="35" place="35" resultid="42151" />
                    <RANKING order="36" place="-1" resultid="43058" />
                    <RANKING order="37" place="-1" resultid="41750" />
                    <RANKING order="38" place="-1" resultid="42100" />
                    <RANKING order="39" place="-1" resultid="43833" />
                    <RANKING order="40" place="-1" resultid="42165" />
                    <RANKING order="41" place="-1" resultid="42024" />
                    <RANKING order="42" place="-1" resultid="42111" />
                    <RANKING order="43" place="-1" resultid="42788" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="44916" daytime="09:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="44917" daytime="09:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="44918" daytime="10:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="44919" daytime="10:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="44920" daytime="10:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="44921" daytime="10:20" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2552" daytime="10:20" gender="F" number="13" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45599" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42501" />
                    <RANKING order="2" place="2" resultid="42994" />
                    <RANKING order="3" place="3" resultid="44029" />
                    <RANKING order="4" place="4" resultid="44034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45600" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41724" />
                    <RANKING order="2" place="2" resultid="43662" />
                    <RANKING order="3" place="3" resultid="43968" />
                    <RANKING order="4" place="4" resultid="42078" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45601" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41994" />
                    <RANKING order="2" place="2" resultid="43557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45602" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="45603" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45604" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43219" />
                    <RANKING order="2" place="2" resultid="41937" />
                    <RANKING order="3" place="3" resultid="43751" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45605" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42135" />
                    <RANKING order="2" place="2" resultid="43757" />
                    <RANKING order="3" place="-1" resultid="41757" />
                    <RANKING order="4" place="-1" resultid="41856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45606" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43850" />
                    <RANKING order="2" place="2" resultid="41745" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45607" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="45608" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="45609" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45610" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45611" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45612" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45613" agemax="-1" agemin="-1" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42501" />
                    <RANKING order="2" place="2" resultid="41724" />
                    <RANKING order="3" place="3" resultid="42994" />
                    <RANKING order="4" place="4" resultid="43662" />
                    <RANKING order="5" place="5" resultid="43968" />
                    <RANKING order="6" place="6" resultid="41994" />
                    <RANKING order="7" place="7" resultid="43219" />
                    <RANKING order="8" place="8" resultid="44029" />
                    <RANKING order="9" place="9" resultid="44034" />
                    <RANKING order="10" place="10" resultid="42078" />
                    <RANKING order="11" place="11" resultid="42135" />
                    <RANKING order="12" place="12" resultid="43251" />
                    <RANKING order="13" place="13" resultid="41937" />
                    <RANKING order="14" place="14" resultid="43557" />
                    <RANKING order="15" place="15" resultid="43757" />
                    <RANKING order="16" place="16" resultid="43751" />
                    <RANKING order="17" place="17" resultid="43850" />
                    <RANKING order="18" place="18" resultid="41745" />
                    <RANKING order="19" place="-1" resultid="41757" />
                    <RANKING order="20" place="-1" resultid="41856" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="44922" daytime="10:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="44923" daytime="10:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="44924" daytime="10:30" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2323" daytime="10:30" gender="M" number="14" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45434" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42702" />
                    <RANKING order="2" place="2" resultid="42325" />
                    <RANKING order="3" place="3" resultid="43934" />
                    <RANKING order="4" place="4" resultid="42819" />
                    <RANKING order="5" place="5" resultid="42375" />
                    <RANKING order="6" place="6" resultid="42866" />
                    <RANKING order="7" place="7" resultid="41733" />
                    <RANKING order="8" place="8" resultid="42676" />
                    <RANKING order="9" place="-1" resultid="42340" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45435" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43743" />
                    <RANKING order="2" place="2" resultid="43892" />
                    <RANKING order="3" place="3" resultid="43148" />
                    <RANKING order="4" place="4" resultid="41978" />
                    <RANKING order="5" place="5" resultid="41950" />
                    <RANKING order="6" place="-1" resultid="41530" />
                    <RANKING order="7" place="-1" resultid="42778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45436" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42484" />
                    <RANKING order="2" place="2" resultid="42766" />
                    <RANKING order="3" place="3" resultid="43918" />
                    <RANKING order="4" place="4" resultid="41876" />
                    <RANKING order="5" place="5" resultid="42033" />
                    <RANKING order="6" place="6" resultid="44852" />
                    <RANKING order="7" place="7" resultid="43719" />
                    <RANKING order="8" place="-1" resultid="42231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45437" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43466" />
                    <RANKING order="2" place="2" resultid="42088" />
                    <RANKING order="3" place="3" resultid="43364" />
                    <RANKING order="4" place="4" resultid="43461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45438" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42198" />
                    <RANKING order="2" place="2" resultid="41791" />
                    <RANKING order="3" place="3" resultid="43548" />
                    <RANKING order="4" place="4" resultid="43448" />
                    <RANKING order="5" place="5" resultid="43723" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45439" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41634" />
                    <RANKING order="2" place="2" resultid="43385" />
                    <RANKING order="3" place="3" resultid="43257" />
                    <RANKING order="4" place="4" resultid="42475" />
                    <RANKING order="5" place="5" resultid="43838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45440" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43803" />
                    <RANKING order="2" place="2" resultid="43071" />
                    <RANKING order="3" place="3" resultid="43191" />
                    <RANKING order="4" place="4" resultid="41671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45441" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="45442" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41694" />
                    <RANKING order="2" place="2" resultid="43020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45443" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42744" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45444" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45445" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45446" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45447" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45448" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43743" />
                    <RANKING order="2" place="2" resultid="42702" />
                    <RANKING order="3" place="3" resultid="42325" />
                    <RANKING order="4" place="4" resultid="43934" />
                    <RANKING order="5" place="5" resultid="42819" />
                    <RANKING order="6" place="6" resultid="42484" />
                    <RANKING order="7" place="7" resultid="43466" />
                    <RANKING order="8" place="8" resultid="42766" />
                    <RANKING order="9" place="9" resultid="42375" />
                    <RANKING order="10" place="10" resultid="43918" />
                    <RANKING order="11" place="11" resultid="41634" />
                    <RANKING order="12" place="12" resultid="43892" />
                    <RANKING order="13" place="13" resultid="42198" />
                    <RANKING order="14" place="14" resultid="42088" />
                    <RANKING order="15" place="15" resultid="43385" />
                    <RANKING order="16" place="16" resultid="41791" />
                    <RANKING order="17" place="17" resultid="41876" />
                    <RANKING order="18" place="18" resultid="42866" />
                    <RANKING order="19" place="19" resultid="41733" />
                    <RANKING order="20" place="20" resultid="43257" />
                    <RANKING order="21" place="21" resultid="43364" />
                    <RANKING order="22" place="22" resultid="42676" />
                    <RANKING order="23" place="23" resultid="41694" />
                    <RANKING order="24" place="24" resultid="42475" />
                    <RANKING order="25" place="25" resultid="43148" />
                    <RANKING order="26" place="26" resultid="41978" />
                    <RANKING order="27" place="27" resultid="41950" />
                    <RANKING order="28" place="28" resultid="43548" />
                    <RANKING order="29" place="29" resultid="43461" />
                    <RANKING order="30" place="30" resultid="43803" />
                    <RANKING order="31" place="31" resultid="42033" />
                    <RANKING order="32" place="32" resultid="44852" />
                    <RANKING order="33" place="33" resultid="43719" />
                    <RANKING order="34" place="34" resultid="43448" />
                    <RANKING order="35" place="35" resultid="43071" />
                    <RANKING order="36" place="36" resultid="43723" />
                    <RANKING order="37" place="37" resultid="43191" />
                    <RANKING order="38" place="38" resultid="42744" />
                    <RANKING order="39" place="39" resultid="43838" />
                    <RANKING order="40" place="40" resultid="43020" />
                    <RANKING order="41" place="41" resultid="41671" />
                    <RANKING order="42" place="-1" resultid="41530" />
                    <RANKING order="43" place="-1" resultid="42231" />
                    <RANKING order="44" place="-1" resultid="42340" />
                    <RANKING order="45" place="-1" resultid="42778" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="44925" daytime="10:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="44926" daytime="10:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="44927" daytime="10:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="44928" daytime="10:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="44929" daytime="10:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="44930" daytime="10:45" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2607" daytime="10:50" gender="F" number="15" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45584" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42331" />
                    <RANKING order="2" place="2" resultid="42357" />
                    <RANKING order="3" place="3" resultid="42847" />
                    <RANKING order="4" place="4" resultid="42738" />
                    <RANKING order="5" place="5" resultid="42185" />
                    <RANKING order="6" place="6" resultid="42361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45585" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43080" />
                    <RANKING order="2" place="2" resultid="43773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45586" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43779" />
                    <RANKING order="2" place="2" resultid="43710" />
                    <RANKING order="3" place="3" resultid="43558" />
                    <RANKING order="4" place="4" resultid="41770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45587" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43063" />
                    <RANKING order="2" place="2" resultid="43896" />
                    <RANKING order="3" place="3" resultid="42732" />
                    <RANKING order="4" place="4" resultid="42506" />
                    <RANKING order="5" place="5" resultid="41547" />
                    <RANKING order="6" place="6" resultid="42162" />
                    <RANKING order="7" place="7" resultid="42850" />
                    <RANKING order="8" place="8" resultid="42725" />
                    <RANKING order="9" place="9" resultid="41621" />
                    <RANKING order="10" place="-1" resultid="42775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45588" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42083" />
                    <RANKING order="2" place="2" resultid="43869" />
                    <RANKING order="3" place="3" resultid="43240" />
                    <RANKING order="4" place="4" resultid="41989" />
                    <RANKING order="5" place="5" resultid="42758" />
                    <RANKING order="6" place="6" resultid="43231" />
                    <RANKING order="7" place="7" resultid="42840" />
                    <RANKING order="8" place="8" resultid="41815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45589" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42459" />
                    <RANKING order="2" place="2" resultid="43301" />
                    <RANKING order="3" place="3" resultid="43752" />
                    <RANKING order="4" place="4" resultid="44013" />
                    <RANKING order="5" place="5" resultid="42242" />
                    <RANKING order="6" place="-1" resultid="43901" />
                    <RANKING order="7" place="-1" resultid="41962" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45590" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42071" />
                    <RANKING order="2" place="2" resultid="43973" />
                    <RANKING order="3" place="3" resultid="42968" />
                    <RANKING order="4" place="4" resultid="43938" />
                    <RANKING order="5" place="5" resultid="43864" />
                    <RANKING order="6" place="6" resultid="43747" />
                    <RANKING order="7" place="7" resultid="42824" />
                    <RANKING order="8" place="8" resultid="42406" />
                    <RANKING order="9" place="9" resultid="42844" />
                    <RANKING order="10" place="-1" resultid="43423" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45591" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41914" />
                    <RANKING order="2" place="2" resultid="41887" />
                    <RANKING order="3" place="3" resultid="43290" />
                    <RANKING order="4" place="4" resultid="42808" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45592" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41690" />
                    <RANKING order="2" place="-1" resultid="43535" />
                    <RANKING order="3" place="-1" resultid="43955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45593" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41819" />
                    <RANKING order="2" place="2" resultid="43226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45594" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45595" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45596" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45597" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45598" agemax="-1" agemin="-1" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43080" />
                    <RANKING order="2" place="2" resultid="42331" />
                    <RANKING order="3" place="3" resultid="43773" />
                    <RANKING order="4" place="4" resultid="42357" />
                    <RANKING order="5" place="5" resultid="42847" />
                    <RANKING order="6" place="6" resultid="42738" />
                    <RANKING order="7" place="7" resultid="42185" />
                    <RANKING order="8" place="8" resultid="43063" />
                    <RANKING order="9" place="9" resultid="43896" />
                    <RANKING order="10" place="10" resultid="42083" />
                    <RANKING order="11" place="11" resultid="42732" />
                    <RANKING order="12" place="12" resultid="43869" />
                    <RANKING order="13" place="13" resultid="42071" />
                    <RANKING order="14" place="14" resultid="42459" />
                    <RANKING order="15" place="15" resultid="42361" />
                    <RANKING order="16" place="16" resultid="43301" />
                    <RANKING order="17" place="17" resultid="41914" />
                    <RANKING order="18" place="18" resultid="43240" />
                    <RANKING order="19" place="19" resultid="42506" />
                    <RANKING order="20" place="20" resultid="41547" />
                    <RANKING order="21" place="21" resultid="42162" />
                    <RANKING order="22" place="22" resultid="43973" />
                    <RANKING order="23" place="23" resultid="41989" />
                    <RANKING order="24" place="24" resultid="43779" />
                    <RANKING order="25" place="25" resultid="42850" />
                    <RANKING order="26" place="26" resultid="42725" />
                    <RANKING order="27" place="27" resultid="42968" />
                    <RANKING order="28" place="28" resultid="43938" />
                    <RANKING order="29" place="29" resultid="42758" />
                    <RANKING order="30" place="30" resultid="43231" />
                    <RANKING order="31" place="31" resultid="43752" />
                    <RANKING order="32" place="32" resultid="44013" />
                    <RANKING order="33" place="33" resultid="43864" />
                    <RANKING order="34" place="34" resultid="41887" />
                    <RANKING order="35" place="35" resultid="42242" />
                    <RANKING order="36" place="36" resultid="43747" />
                    <RANKING order="37" place="37" resultid="42840" />
                    <RANKING order="38" place="38" resultid="43710" />
                    <RANKING order="39" place="39" resultid="42824" />
                    <RANKING order="40" place="40" resultid="41621" />
                    <RANKING order="41" place="41" resultid="43290" />
                    <RANKING order="42" place="42" resultid="42406" />
                    <RANKING order="43" place="43" resultid="43558" />
                    <RANKING order="44" place="44" resultid="41690" />
                    <RANKING order="45" place="45" resultid="42844" />
                    <RANKING order="46" place="46" resultid="41815" />
                    <RANKING order="47" place="47" resultid="41770" />
                    <RANKING order="48" place="48" resultid="42808" />
                    <RANKING order="49" place="49" resultid="41819" />
                    <RANKING order="50" place="50" resultid="43226" />
                    <RANKING order="51" place="-1" resultid="42775" />
                    <RANKING order="52" place="-1" resultid="43423" />
                    <RANKING order="53" place="-1" resultid="43535" />
                    <RANKING order="54" place="-1" resultid="43901" />
                    <RANKING order="55" place="-1" resultid="43955" />
                    <RANKING order="56" place="-1" resultid="41962" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45097" daytime="10:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45098" daytime="10:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="45099" daytime="10:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="45100" daytime="10:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="45101" daytime="11:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="45102" daytime="11:00" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="45103" daytime="11:05" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2188" daytime="11:05" gender="M" number="16" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45419" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42669" />
                    <RANKING order="2" place="2" resultid="42796" />
                    <RANKING order="3" place="3" resultid="42685" />
                    <RANKING order="4" place="4" resultid="43084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45420" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43930" />
                    <RANKING order="2" place="2" resultid="43685" />
                    <RANKING order="3" place="3" resultid="42710" />
                    <RANKING order="4" place="4" resultid="43134" />
                    <RANKING order="5" place="5" resultid="42432" />
                    <RANKING order="6" place="6" resultid="41985" />
                    <RANKING order="7" place="7" resultid="43784" />
                    <RANKING order="8" place="8" resultid="43162" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45421" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42232" />
                    <RANKING order="2" place="2" resultid="43812" />
                    <RANKING order="3" place="3" resultid="43807" />
                    <RANKING order="4" place="4" resultid="41981" />
                    <RANKING order="5" place="5" resultid="44007" />
                    <RANKING order="6" place="6" resultid="42054" />
                    <RANKING order="7" place="7" resultid="43167" />
                    <RANKING order="8" place="8" resultid="43793" />
                    <RANKING order="9" place="9" resultid="42448" />
                    <RANKING order="10" place="10" resultid="41802" />
                    <RANKING order="11" place="-1" resultid="43089" />
                    <RANKING order="12" place="-1" resultid="43143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45422" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42470" />
                    <RANKING order="2" place="2" resultid="44020" />
                    <RANKING order="3" place="3" resultid="42190" />
                    <RANKING order="4" place="4" resultid="44002" />
                    <RANKING order="5" place="5" resultid="43687" />
                    <RANKING order="6" place="6" resultid="41837" />
                    <RANKING order="7" place="7" resultid="43714" />
                    <RANKING order="8" place="8" resultid="43733" />
                    <RANKING order="9" place="9" resultid="43979" />
                    <RANKING order="10" place="10" resultid="42858" />
                    <RANKING order="11" place="11" resultid="41833" />
                    <RANKING order="12" place="12" resultid="42801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45423" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43587" />
                    <RANKING order="2" place="2" resultid="41845" />
                    <RANKING order="3" place="3" resultid="42962" />
                    <RANKING order="4" place="4" resultid="41809" />
                    <RANKING order="5" place="5" resultid="43598" />
                    <RANKING order="6" place="6" resultid="41867" />
                    <RANKING order="7" place="7" resultid="43910" />
                    <RANKING order="8" place="8" resultid="43990" />
                    <RANKING order="9" place="9" resultid="42417" />
                    <RANKING order="10" place="-1" resultid="43031" />
                    <RANKING order="11" place="-1" resultid="41618" />
                    <RANKING order="12" place="-1" resultid="43442" />
                    <RANKING order="13" place="-1" resultid="43628" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45424" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42489" />
                    <RANKING order="2" place="2" resultid="41899" />
                    <RANKING order="3" place="3" resultid="43282" />
                    <RANKING order="4" place="4" resultid="42984" />
                    <RANKING order="5" place="5" resultid="42213" />
                    <RANKING order="6" place="6" resultid="41629" />
                    <RANKING order="7" place="7" resultid="43763" />
                    <RANKING order="8" place="8" resultid="43591" />
                    <RANKING order="9" place="9" resultid="43185" />
                    <RANKING order="10" place="10" resultid="42862" />
                    <RANKING order="11" place="11" resultid="43157" />
                    <RANKING order="12" place="12" resultid="43728" />
                    <RANKING order="13" place="13" resultid="42411" />
                    <RANKING order="14" place="14" resultid="43051" />
                    <RANKING order="15" place="-1" resultid="42791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45425" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43564" />
                    <RANKING order="2" place="2" resultid="43206" />
                    <RANKING order="3" place="3" resultid="41717" />
                    <RANKING order="4" place="4" resultid="43620" />
                    <RANKING order="5" place="5" resultid="41894" />
                    <RANKING order="6" place="6" resultid="42364" />
                    <RANKING order="7" place="7" resultid="42145" />
                    <RANKING order="8" place="8" resultid="42000" />
                    <RANKING order="9" place="9" resultid="43576" />
                    <RANKING order="10" place="10" resultid="43016" />
                    <RANKING order="11" place="11" resultid="42438" />
                    <RANKING order="12" place="12" resultid="42166" />
                    <RANKING order="13" place="-1" resultid="43964" />
                    <RANKING order="14" place="-1" resultid="42755" />
                    <RANKING order="15" place="-1" resultid="42979" />
                    <RANKING order="16" place="-1" resultid="43509" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45426" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43215" />
                    <RANKING order="2" place="2" resultid="42127" />
                    <RANKING order="3" place="-1" resultid="43514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45427" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41695" />
                    <RANKING order="2" place="2" resultid="42101" />
                    <RANKING order="3" place="3" resultid="43265" />
                    <RANKING order="4" place="4" resultid="41763" />
                    <RANKING order="5" place="5" resultid="41700" />
                    <RANKING order="6" place="6" resultid="42750" />
                    <RANKING order="7" place="7" resultid="42494" />
                    <RANKING order="8" place="8" resultid="43391" />
                    <RANKING order="9" place="9" resultid="43153" />
                    <RANKING order="10" place="10" resultid="42152" />
                    <RANKING order="11" place="11" resultid="43495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45428" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41871" />
                    <RANKING order="2" place="2" resultid="42414" />
                    <RANKING order="3" place="3" resultid="43359" />
                    <RANKING order="4" place="4" resultid="41677" />
                    <RANKING order="5" place="5" resultid="42403" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45429" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41665" />
                    <RANKING order="2" place="2" resultid="43541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45430" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45431" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45432" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45433" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43930" />
                    <RANKING order="2" place="2" resultid="43587" />
                    <RANKING order="3" place="3" resultid="43685" />
                    <RANKING order="4" place="4" resultid="42669" />
                    <RANKING order="5" place="5" resultid="41845" />
                    <RANKING order="6" place="6" resultid="42796" />
                    <RANKING order="7" place="7" resultid="42470" />
                    <RANKING order="8" place="8" resultid="42232" />
                    <RANKING order="9" place="9" resultid="42710" />
                    <RANKING order="10" place="10" resultid="43134" />
                    <RANKING order="11" place="11" resultid="43812" />
                    <RANKING order="12" place="12" resultid="43564" />
                    <RANKING order="13" place="13" resultid="43807" />
                    <RANKING order="14" place="14" resultid="43206" />
                    <RANKING order="15" place="15" resultid="42685" />
                    <RANKING order="16" place="16" resultid="44020" />
                    <RANKING order="17" place="17" resultid="42489" />
                    <RANKING order="18" place="18" resultid="42190" />
                    <RANKING order="19" place="19" resultid="41899" />
                    <RANKING order="20" place="20" resultid="43282" />
                    <RANKING order="21" place="21" resultid="43215" />
                    <RANKING order="22" place="22" resultid="42432" />
                    <RANKING order="23" place="23" resultid="43084" />
                    <RANKING order="24" place="24" resultid="42984" />
                    <RANKING order="25" place="25" resultid="41981" />
                    <RANKING order="26" place="26" resultid="41985" />
                    <RANKING order="27" place="27" resultid="42962" />
                    <RANKING order="28" place="28" resultid="44007" />
                    <RANKING order="29" place="29" resultid="43784" />
                    <RANKING order="30" place="30" resultid="42054" />
                    <RANKING order="31" place="31" resultid="44002" />
                    <RANKING order="32" place="32" resultid="41809" />
                    <RANKING order="33" place="33" resultid="43598" />
                    <RANKING order="34" place="34" resultid="41717" />
                    <RANKING order="35" place="35" resultid="42213" />
                    <RANKING order="36" place="36" resultid="43167" />
                    <RANKING order="37" place="37" resultid="43687" />
                    <RANKING order="38" place="38" resultid="41867" />
                    <RANKING order="39" place="39" resultid="41837" />
                    <RANKING order="40" place="40" resultid="43714" />
                    <RANKING order="41" place="41" resultid="43910" />
                    <RANKING order="42" place="42" resultid="41629" />
                    <RANKING order="43" place="43" resultid="43620" />
                    <RANKING order="44" place="44" resultid="41894" />
                    <RANKING order="45" place="45" resultid="43990" />
                    <RANKING order="46" place="46" resultid="42364" />
                    <RANKING order="47" place="47" resultid="42417" />
                    <RANKING order="48" place="48" resultid="41695" />
                    <RANKING order="49" place="48" resultid="43763" />
                    <RANKING order="50" place="50" resultid="43591" />
                    <RANKING order="51" place="51" resultid="42101" />
                    <RANKING order="52" place="52" resultid="42145" />
                    <RANKING order="53" place="52" resultid="43185" />
                    <RANKING order="54" place="54" resultid="43793" />
                    <RANKING order="55" place="55" resultid="42000" />
                    <RANKING order="56" place="56" resultid="43576" />
                    <RANKING order="57" place="57" resultid="43162" />
                    <RANKING order="58" place="58" resultid="41871" />
                    <RANKING order="59" place="59" resultid="43733" />
                    <RANKING order="60" place="60" resultid="43016" />
                    <RANKING order="61" place="61" resultid="43979" />
                    <RANKING order="62" place="62" resultid="42862" />
                    <RANKING order="63" place="63" resultid="42858" />
                    <RANKING order="64" place="64" resultid="43265" />
                    <RANKING order="65" place="65" resultid="43157" />
                    <RANKING order="66" place="66" resultid="41833" />
                    <RANKING order="67" place="67" resultid="41763" />
                    <RANKING order="68" place="68" resultid="42801" />
                    <RANKING order="69" place="69" resultid="43728" />
                    <RANKING order="70" place="70" resultid="41700" />
                    <RANKING order="71" place="71" resultid="42448" />
                    <RANKING order="72" place="72" resultid="42414" />
                    <RANKING order="73" place="73" resultid="41665" />
                    <RANKING order="74" place="74" resultid="42750" />
                    <RANKING order="75" place="75" resultid="42494" />
                    <RANKING order="76" place="76" resultid="42411" />
                    <RANKING order="77" place="77" resultid="42438" />
                    <RANKING order="78" place="78" resultid="41802" />
                    <RANKING order="79" place="79" resultid="43391" />
                    <RANKING order="80" place="80" resultid="43541" />
                    <RANKING order="81" place="81" resultid="43153" />
                    <RANKING order="82" place="82" resultid="43051" />
                    <RANKING order="83" place="83" resultid="43359" />
                    <RANKING order="84" place="84" resultid="42152" />
                    <RANKING order="85" place="85" resultid="42166" />
                    <RANKING order="86" place="86" resultid="43495" />
                    <RANKING order="87" place="87" resultid="41677" />
                    <RANKING order="88" place="88" resultid="42403" />
                    <RANKING order="89" place="89" resultid="41905" />
                    <RANKING order="90" place="90" resultid="42127" />
                    <RANKING order="91" place="-1" resultid="43089" />
                    <RANKING order="92" place="-1" resultid="43964" />
                    <RANKING order="93" place="-1" resultid="43031" />
                    <RANKING order="94" place="-1" resultid="41618" />
                    <RANKING order="95" place="-1" resultid="42755" />
                    <RANKING order="96" place="-1" resultid="42791" />
                    <RANKING order="97" place="-1" resultid="42979" />
                    <RANKING order="98" place="-1" resultid="43143" />
                    <RANKING order="99" place="-1" resultid="43442" />
                    <RANKING order="100" place="-1" resultid="43509" />
                    <RANKING order="101" place="-1" resultid="43514" />
                    <RANKING order="102" place="-1" resultid="43628" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="44938" daytime="11:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="44939" daytime="11:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="44940" daytime="11:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="44941" daytime="11:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="44942" daytime="11:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="44943" daytime="11:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="44944" daytime="11:20" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="44945" daytime="11:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="44946" daytime="11:20" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="44947" daytime="11:25" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="44948" daytime="11:25" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="44949" daytime="11:30" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="44950" daytime="11:30" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2021-07-10" daytime="15:00" endtime="17:11" name="2ª Jornada-2ª sessão" number="4">
          <EVENTS>
            <EVENT eventid="2637" daytime="15:00" gender="F" number="17" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45569" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42332" />
                    <RANKING order="2" place="2" resultid="43668" />
                    <RANKING order="3" place="3" resultid="42454" />
                    <RANKING order="4" place="4" resultid="42995" />
                    <RANKING order="5" place="5" resultid="42352" />
                    <RANKING order="6" place="6" resultid="42158" />
                    <RANKING order="7" place="7" resultid="42464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45570" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43774" />
                    <RANKING order="2" place="2" resultid="42202" />
                    <RANKING order="3" place="3" resultid="42079" />
                    <RANKING order="4" place="4" resultid="43637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45571" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43412" />
                    <RANKING order="2" place="2" resultid="42237" />
                    <RANKING order="3" place="3" resultid="43559" />
                    <RANKING order="4" place="-1" resultid="41525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45572" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43064" />
                    <RANKING order="2" place="2" resultid="43039" />
                    <RANKING order="3" place="3" resultid="43906" />
                    <RANKING order="4" place="4" resultid="42507" />
                    <RANKING order="5" place="5" resultid="41548" />
                    <RANKING order="6" place="6" resultid="42851" />
                    <RANKING order="7" place="7" resultid="41622" />
                    <RANKING order="8" place="-1" resultid="42776" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45573" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42084" />
                    <RANKING order="2" place="2" resultid="41972" />
                    <RANKING order="3" place="3" resultid="42759" />
                    <RANKING order="4" place="4" resultid="41945" />
                    <RANKING order="5" place="5" resultid="42715" />
                    <RANKING order="6" place="6" resultid="42841" />
                    <RANKING order="7" place="-1" resultid="41941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45574" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43302" />
                    <RANKING order="2" place="2" resultid="44014" />
                    <RANKING order="3" place="3" resultid="43902" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45575" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42140" />
                    <RANKING order="2" place="2" resultid="43331" />
                    <RANKING order="3" place="3" resultid="43974" />
                    <RANKING order="4" place="4" resultid="41920" />
                    <RANKING order="5" place="5" resultid="43865" />
                    <RANKING order="6" place="6" resultid="43758" />
                    <RANKING order="7" place="7" resultid="42691" />
                    <RANKING order="8" place="8" resultid="41758" />
                    <RANKING order="9" place="9" resultid="43478" />
                    <RANKING order="10" place="10" resultid="43651" />
                    <RANKING order="11" place="11" resultid="42845" />
                    <RANKING order="12" place="-1" resultid="43424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45576" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41915" />
                    <RANKING order="2" place="2" resultid="43851" />
                    <RANKING order="3" place="3" resultid="43644" />
                    <RANKING order="4" place="4" resultid="43139" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45577" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41882" />
                    <RANKING order="2" place="2" resultid="41691" />
                    <RANKING order="3" place="3" resultid="43536" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45578" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43227" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45579" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45580" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45581" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45582" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45583" agemax="-1" agemin="-1" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42332" />
                    <RANKING order="2" place="2" resultid="43668" />
                    <RANKING order="3" place="3" resultid="42454" />
                    <RANKING order="4" place="4" resultid="42995" />
                    <RANKING order="5" place="5" resultid="42084" />
                    <RANKING order="6" place="6" resultid="43412" />
                    <RANKING order="7" place="7" resultid="43774" />
                    <RANKING order="8" place="8" resultid="43064" />
                    <RANKING order="9" place="9" resultid="42352" />
                    <RANKING order="10" place="10" resultid="42202" />
                    <RANKING order="11" place="11" resultid="43302" />
                    <RANKING order="12" place="12" resultid="42140" />
                    <RANKING order="13" place="13" resultid="43039" />
                    <RANKING order="14" place="14" resultid="43906" />
                    <RANKING order="15" place="15" resultid="42158" />
                    <RANKING order="16" place="16" resultid="41972" />
                    <RANKING order="17" place="17" resultid="42079" />
                    <RANKING order="18" place="18" resultid="43637" />
                    <RANKING order="19" place="19" resultid="42464" />
                    <RANKING order="20" place="20" resultid="42507" />
                    <RANKING order="21" place="21" resultid="43331" />
                    <RANKING order="22" place="22" resultid="43974" />
                    <RANKING order="23" place="23" resultid="41920" />
                    <RANKING order="24" place="24" resultid="42759" />
                    <RANKING order="25" place="25" resultid="41915" />
                    <RANKING order="26" place="26" resultid="43865" />
                    <RANKING order="27" place="27" resultid="41945" />
                    <RANKING order="28" place="28" resultid="41548" />
                    <RANKING order="29" place="29" resultid="42851" />
                    <RANKING order="30" place="30" resultid="42715" />
                    <RANKING order="31" place="30" resultid="43851" />
                    <RANKING order="32" place="32" resultid="42237" />
                    <RANKING order="33" place="33" resultid="42841" />
                    <RANKING order="34" place="34" resultid="43758" />
                    <RANKING order="35" place="35" resultid="43559" />
                    <RANKING order="36" place="36" resultid="42691" />
                    <RANKING order="37" place="37" resultid="44014" />
                    <RANKING order="38" place="38" resultid="41758" />
                    <RANKING order="39" place="39" resultid="41882" />
                    <RANKING order="40" place="40" resultid="43902" />
                    <RANKING order="41" place="41" resultid="41622" />
                    <RANKING order="42" place="42" resultid="43478" />
                    <RANKING order="43" place="43" resultid="43651" />
                    <RANKING order="44" place="44" resultid="43644" />
                    <RANKING order="45" place="45" resultid="41691" />
                    <RANKING order="46" place="46" resultid="42845" />
                    <RANKING order="47" place="47" resultid="43536" />
                    <RANKING order="48" place="48" resultid="43139" />
                    <RANKING order="49" place="49" resultid="43227" />
                    <RANKING order="50" place="-1" resultid="42776" />
                    <RANKING order="51" place="-1" resultid="43424" />
                    <RANKING order="52" place="-1" resultid="41525" />
                    <RANKING order="53" place="-1" resultid="41941" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="44951" daytime="15:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="44952" daytime="15:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="44953" daytime="15:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="44954" daytime="15:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="44955" daytime="15:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="44956" daytime="15:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="44957" daytime="15:20" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2415" daytime="15:20" gender="M" number="18" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45404" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41824" />
                    <RANKING order="2" place="2" resultid="42326" />
                    <RANKING order="3" place="3" resultid="42703" />
                    <RANKING order="4" place="4" resultid="42820" />
                    <RANKING order="5" place="5" resultid="43935" />
                    <RANKING order="6" place="6" resultid="42797" />
                    <RANKING order="7" place="7" resultid="42370" />
                    <RANKING order="8" place="8" resultid="42835" />
                    <RANKING order="9" place="9" resultid="41734" />
                    <RANKING order="10" place="10" resultid="42686" />
                    <RANKING order="11" place="11" resultid="42867" />
                    <RANKING order="12" place="12" resultid="43704" />
                    <RANKING order="13" place="-1" resultid="42341" />
                    <RANKING order="14" place="-1" resultid="42814" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45405" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42105" />
                    <RANKING order="2" place="2" resultid="43744" />
                    <RANKING order="3" place="3" resultid="42433" />
                    <RANKING order="4" place="4" resultid="43674" />
                    <RANKING order="5" place="5" resultid="43306" />
                    <RANKING order="6" place="6" resultid="43149" />
                    <RANKING order="7" place="7" resultid="43654" />
                    <RANKING order="8" place="8" resultid="43632" />
                    <RANKING order="9" place="9" resultid="41986" />
                    <RANKING order="10" place="10" resultid="41979" />
                    <RANKING order="11" place="11" resultid="43785" />
                    <RANKING order="12" place="12" resultid="43163" />
                    <RANKING order="13" place="13" resultid="41951" />
                    <RANKING order="14" place="-1" resultid="41531" />
                    <RANKING order="15" place="-1" resultid="42025" />
                    <RANKING order="16" place="-1" resultid="43860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45406" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42772" />
                    <RANKING order="2" place="2" resultid="43473" />
                    <RANKING order="3" place="3" resultid="42485" />
                    <RANKING order="4" place="4" resultid="41982" />
                    <RANKING order="5" place="5" resultid="43813" />
                    <RANKING order="6" place="6" resultid="43700" />
                    <RANKING order="7" place="7" resultid="42767" />
                    <RANKING order="8" place="8" resultid="43168" />
                    <RANKING order="9" place="9" resultid="43720" />
                    <RANKING order="10" place="10" resultid="41647" />
                    <RANKING order="11" place="11" resultid="42449" />
                    <RANKING order="12" place="12" resultid="44853" />
                    <RANKING order="13" place="13" resultid="41803" />
                    <RANKING order="14" place="-1" resultid="43144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45407" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43467" />
                    <RANKING order="2" place="2" resultid="41924" />
                    <RANKING order="3" place="3" resultid="43795" />
                    <RANKING order="4" place="4" resultid="43462" />
                    <RANKING order="5" place="5" resultid="41838" />
                    <RANKING order="6" place="6" resultid="42247" />
                    <RANKING order="7" place="7" resultid="42802" />
                    <RANKING order="8" place="-1" resultid="43403" />
                    <RANKING order="9" place="-1" resultid="41520" />
                    <RANKING order="10" place="-1" resultid="41957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45408" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43175" />
                    <RANKING order="2" place="2" resultid="43549" />
                    <RANKING order="3" place="3" resultid="42963" />
                    <RANKING order="4" place="4" resultid="43378" />
                    <RANKING order="5" place="5" resultid="42956" />
                    <RANKING order="6" place="6" resultid="42429" />
                    <RANKING order="7" place="7" resultid="43991" />
                    <RANKING order="8" place="8" resultid="43420" />
                    <RANKING order="9" place="9" resultid="41738" />
                    <RANKING order="10" place="10" resultid="43724" />
                    <RANKING order="11" place="11" resultid="43911" />
                    <RANKING order="12" place="12" resultid="43032" />
                    <RANKING order="13" place="-1" resultid="41795" />
                    <RANKING order="14" place="-1" resultid="43855" />
                    <RANKING order="15" place="-1" resultid="43986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45409" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43386" />
                    <RANKING order="2" place="2" resultid="42219" />
                    <RANKING order="3" place="3" resultid="43258" />
                    <RANKING order="4" place="4" resultid="43283" />
                    <RANKING order="5" place="5" resultid="43887" />
                    <RANKING order="6" place="6" resultid="41627" />
                    <RANKING order="7" place="7" resultid="43592" />
                    <RANKING order="8" place="8" resultid="44025" />
                    <RANKING order="9" place="9" resultid="43186" />
                    <RANKING order="10" place="10" resultid="43834" />
                    <RANKING order="11" place="11" resultid="43351" />
                    <RANKING order="12" place="12" resultid="43729" />
                    <RANKING order="13" place="13" resultid="43158" />
                    <RANKING order="14" place="-1" resultid="43505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45410" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43612" />
                    <RANKING order="2" place="2" resultid="41718" />
                    <RANKING order="3" place="3" resultid="43192" />
                    <RANKING order="4" place="4" resultid="42146" />
                    <RANKING order="5" place="5" resultid="42365" />
                    <RANKING order="6" place="-1" resultid="43577" />
                    <RANKING order="7" place="-1" resultid="43925" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45411" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41686" />
                    <RANKING order="2" place="2" resultid="43515" />
                    <RANKING order="3" place="3" resultid="42116" />
                    <RANKING order="4" place="4" resultid="42039" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45412" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41696" />
                    <RANKING order="2" place="2" resultid="41764" />
                    <RANKING order="3" place="3" resultid="42751" />
                    <RANKING order="4" place="4" resultid="43392" />
                    <RANKING order="5" place="5" resultid="43021" />
                    <RANKING order="6" place="6" resultid="43027" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45413" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45414" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45415" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45416" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45417" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45418" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42105" />
                    <RANKING order="2" place="2" resultid="41824" />
                    <RANKING order="3" place="3" resultid="42326" />
                    <RANKING order="4" place="4" resultid="42703" />
                    <RANKING order="5" place="5" resultid="42772" />
                    <RANKING order="6" place="6" resultid="42820" />
                    <RANKING order="7" place="7" resultid="43744" />
                    <RANKING order="8" place="8" resultid="43473" />
                    <RANKING order="9" place="9" resultid="43935" />
                    <RANKING order="10" place="10" resultid="42797" />
                    <RANKING order="11" place="11" resultid="42485" />
                    <RANKING order="12" place="12" resultid="43175" />
                    <RANKING order="13" place="13" resultid="43386" />
                    <RANKING order="14" place="14" resultid="43467" />
                    <RANKING order="15" place="15" resultid="42370" />
                    <RANKING order="16" place="16" resultid="42835" />
                    <RANKING order="17" place="17" resultid="43612" />
                    <RANKING order="18" place="18" resultid="42433" />
                    <RANKING order="19" place="19" resultid="43674" />
                    <RANKING order="20" place="20" resultid="42219" />
                    <RANKING order="21" place="21" resultid="43306" />
                    <RANKING order="22" place="22" resultid="41982" />
                    <RANKING order="23" place="23" resultid="43813" />
                    <RANKING order="24" place="24" resultid="41924" />
                    <RANKING order="25" place="25" resultid="43549" />
                    <RANKING order="26" place="26" resultid="43700" />
                    <RANKING order="27" place="27" resultid="43149" />
                    <RANKING order="28" place="28" resultid="42767" />
                    <RANKING order="29" place="29" resultid="41734" />
                    <RANKING order="30" place="30" resultid="43258" />
                    <RANKING order="31" place="31" resultid="43654" />
                    <RANKING order="32" place="32" resultid="42686" />
                    <RANKING order="33" place="33" resultid="43632" />
                    <RANKING order="34" place="34" resultid="41986" />
                    <RANKING order="35" place="35" resultid="43283" />
                    <RANKING order="36" place="36" resultid="41686" />
                    <RANKING order="37" place="37" resultid="41979" />
                    <RANKING order="38" place="38" resultid="41696" />
                    <RANKING order="39" place="39" resultid="41718" />
                    <RANKING order="40" place="40" resultid="43785" />
                    <RANKING order="41" place="41" resultid="42867" />
                    <RANKING order="42" place="42" resultid="42963" />
                    <RANKING order="43" place="43" resultid="43887" />
                    <RANKING order="44" place="44" resultid="43795" />
                    <RANKING order="45" place="45" resultid="43704" />
                    <RANKING order="46" place="46" resultid="43378" />
                    <RANKING order="47" place="47" resultid="43515" />
                    <RANKING order="48" place="48" resultid="43462" />
                    <RANKING order="49" place="49" resultid="43163" />
                    <RANKING order="50" place="50" resultid="43168" />
                    <RANKING order="51" place="51" resultid="41838" />
                    <RANKING order="52" place="52" resultid="42956" />
                    <RANKING order="53" place="53" resultid="43720" />
                    <RANKING order="54" place="54" resultid="42247" />
                    <RANKING order="55" place="55" resultid="42429" />
                    <RANKING order="56" place="56" resultid="41627" />
                    <RANKING order="57" place="57" resultid="42116" />
                    <RANKING order="58" place="58" resultid="43991" />
                    <RANKING order="59" place="59" resultid="41951" />
                    <RANKING order="60" place="60" resultid="43420" />
                    <RANKING order="61" place="61" resultid="41661" />
                    <RANKING order="62" place="62" resultid="41647" />
                    <RANKING order="63" place="63" resultid="41738" />
                    <RANKING order="64" place="64" resultid="43724" />
                    <RANKING order="65" place="65" resultid="43592" />
                    <RANKING order="66" place="66" resultid="42449" />
                    <RANKING order="67" place="67" resultid="44025" />
                    <RANKING order="68" place="68" resultid="43192" />
                    <RANKING order="69" place="69" resultid="44853" />
                    <RANKING order="70" place="70" resultid="43911" />
                    <RANKING order="71" place="71" resultid="42146" />
                    <RANKING order="72" place="72" resultid="41764" />
                    <RANKING order="73" place="73" resultid="42365" />
                    <RANKING order="74" place="74" resultid="43186" />
                    <RANKING order="75" place="75" resultid="43834" />
                    <RANKING order="76" place="76" resultid="43032" />
                    <RANKING order="77" place="77" resultid="42039" />
                    <RANKING order="78" place="78" resultid="43351" />
                    <RANKING order="79" place="79" resultid="42802" />
                    <RANKING order="80" place="80" resultid="42751" />
                    <RANKING order="81" place="81" resultid="43729" />
                    <RANKING order="82" place="82" resultid="43392" />
                    <RANKING order="83" place="83" resultid="41654" />
                    <RANKING order="84" place="84" resultid="43158" />
                    <RANKING order="85" place="85" resultid="43021" />
                    <RANKING order="86" place="86" resultid="43027" />
                    <RANKING order="87" place="87" resultid="41803" />
                    <RANKING order="88" place="-1" resultid="43505" />
                    <RANKING order="89" place="-1" resultid="41531" />
                    <RANKING order="90" place="-1" resultid="41795" />
                    <RANKING order="91" place="-1" resultid="42025" />
                    <RANKING order="92" place="-1" resultid="42341" />
                    <RANKING order="93" place="-1" resultid="42814" />
                    <RANKING order="94" place="-1" resultid="43144" />
                    <RANKING order="95" place="-1" resultid="43403" />
                    <RANKING order="96" place="-1" resultid="43577" />
                    <RANKING order="97" place="-1" resultid="43855" />
                    <RANKING order="98" place="-1" resultid="43860" />
                    <RANKING order="99" place="-1" resultid="43925" />
                    <RANKING order="100" place="-1" resultid="41520" />
                    <RANKING order="101" place="-1" resultid="41957" />
                    <RANKING order="102" place="-1" resultid="43986" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45104" daytime="15:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45105" daytime="15:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="45106" daytime="15:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="45107" daytime="15:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="45108" daytime="15:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="45109" daytime="15:35" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="45110" daytime="15:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="45111" daytime="15:40" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="45112" daytime="15:45" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="45113" daytime="15:45" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="45114" daytime="15:50" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="45115" daytime="15:50" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="45116" daytime="15:55" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2233" daytime="15:55" gender="F" number="19" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45554" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42502" />
                    <RANKING order="2" place="2" resultid="43960" />
                    <RANKING order="3" place="3" resultid="44035" />
                    <RANKING order="4" place="4" resultid="44030" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45555" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43969" />
                    <RANKING order="2" place="2" resultid="42443" />
                    <RANKING order="3" place="3" resultid="43641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45556" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42421" />
                    <RANKING order="2" place="2" resultid="43413" />
                    <RANKING order="3" place="3" resultid="43560" />
                    <RANKING order="4" place="-1" resultid="41771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45557" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43065" />
                    <RANKING order="2" place="2" resultid="42697" />
                    <RANKING order="3" place="3" resultid="43897" />
                    <RANKING order="4" place="4" resultid="43040" />
                    <RANKING order="5" place="5" resultid="43047" />
                    <RANKING order="6" place="-1" resultid="43528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45558" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42121" />
                    <RANKING order="2" place="2" resultid="43279" />
                    <RANKING order="3" place="3" resultid="43870" />
                    <RANKING order="4" place="4" resultid="43241" />
                    <RANKING order="5" place="5" resultid="43252" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45559" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42046" />
                    <RANKING order="2" place="2" resultid="42175" />
                    <RANKING order="3" place="3" resultid="43680" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45560" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41921" />
                    <RANKING order="2" place="2" resultid="43125" />
                    <RANKING order="3" place="3" resultid="43479" />
                    <RANKING order="4" place="-1" resultid="43373" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45561" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41746" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45562" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="45563" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="45564" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45565" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45566" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45567" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45568" agemax="-1" agemin="-1" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42502" />
                    <RANKING order="2" place="2" resultid="43960" />
                    <RANKING order="3" place="3" resultid="42121" />
                    <RANKING order="4" place="4" resultid="43969" />
                    <RANKING order="5" place="5" resultid="42421" />
                    <RANKING order="6" place="6" resultid="43279" />
                    <RANKING order="7" place="7" resultid="43065" />
                    <RANKING order="8" place="8" resultid="42046" />
                    <RANKING order="9" place="9" resultid="42697" />
                    <RANKING order="10" place="10" resultid="43413" />
                    <RANKING order="11" place="11" resultid="43870" />
                    <RANKING order="12" place="12" resultid="44035" />
                    <RANKING order="13" place="13" resultid="43897" />
                    <RANKING order="14" place="14" resultid="42443" />
                    <RANKING order="15" place="15" resultid="44030" />
                    <RANKING order="16" place="16" resultid="43040" />
                    <RANKING order="17" place="17" resultid="43241" />
                    <RANKING order="18" place="18" resultid="43641" />
                    <RANKING order="19" place="19" resultid="41921" />
                    <RANKING order="20" place="20" resultid="43252" />
                    <RANKING order="21" place="21" resultid="42175" />
                    <RANKING order="22" place="22" resultid="43047" />
                    <RANKING order="23" place="23" resultid="43560" />
                    <RANKING order="24" place="24" resultid="43680" />
                    <RANKING order="25" place="25" resultid="43125" />
                    <RANKING order="26" place="26" resultid="41746" />
                    <RANKING order="27" place="27" resultid="43479" />
                    <RANKING order="28" place="-1" resultid="41771" />
                    <RANKING order="29" place="-1" resultid="43373" />
                    <RANKING order="30" place="-1" resultid="43528" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="44971" daytime="15:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="44972" daytime="16:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="44973" daytime="16:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="44974" daytime="16:15" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2385" daytime="16:15" gender="M" number="20" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45389" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42821" />
                    <RANKING order="2" place="2" resultid="43085" />
                    <RANKING order="3" place="3" resultid="42868" />
                    <RANKING order="4" place="4" resultid="42677" />
                    <RANKING order="5" place="-1" resultid="43738" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45390" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42779" />
                    <RANKING order="2" place="2" resultid="43893" />
                    <RANKING order="3" place="3" resultid="42012" />
                    <RANKING order="4" place="4" resultid="43307" />
                    <RANKING order="5" place="5" resultid="43135" />
                    <RANKING order="6" place="6" resultid="43675" />
                    <RANKING order="7" place="7" resultid="42019" />
                    <RANKING order="8" place="-1" resultid="43150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45391" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43822" />
                    <RANKING order="2" place="2" resultid="43946" />
                    <RANKING order="3" place="3" resultid="42050" />
                    <RANKING order="4" place="4" resultid="43919" />
                    <RANKING order="5" place="5" resultid="41877" />
                    <RANKING order="6" place="6" resultid="44008" />
                    <RANKING order="7" place="7" resultid="41983" />
                    <RANKING order="8" place="8" resultid="43076" />
                    <RANKING order="9" place="9" resultid="44854" />
                    <RANKING order="10" place="10" resultid="43409" />
                    <RANKING order="11" place="-1" resultid="42061" />
                    <RANKING order="12" place="-1" resultid="41830" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45392" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42989" />
                    <RANKING order="2" place="2" resultid="43943" />
                    <RANKING order="3" place="3" resultid="43365" />
                    <RANKING order="4" place="4" resultid="41910" />
                    <RANKING order="5" place="5" resultid="42191" />
                    <RANKING order="6" place="6" resultid="43463" />
                    <RANKING order="7" place="7" resultid="41834" />
                    <RANKING order="8" place="8" resultid="41751" />
                    <RANKING order="9" place="9" resultid="43980" />
                    <RANKING order="10" place="10" resultid="43696" />
                    <RANKING order="11" place="-1" resultid="44003" />
                    <RANKING order="12" place="-1" resultid="42066" />
                    <RANKING order="13" place="-1" resultid="43468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45393" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41810" />
                    <RANKING order="2" place="2" resultid="41967" />
                    <RANKING order="3" place="3" resultid="41739" />
                    <RANKING order="4" place="4" resultid="43532" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45394" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42476" />
                    <RANKING order="2" place="2" resultid="41900" />
                    <RANKING order="3" place="3" resultid="42181" />
                    <RANKING order="4" place="4" resultid="43888" />
                    <RANKING order="5" place="5" resultid="43839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45395" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43346" />
                    <RANKING order="2" place="2" resultid="41719" />
                    <RANKING order="3" place="3" resultid="42001" />
                    <RANKING order="4" place="4" resultid="41860" />
                    <RANKING order="5" place="5" resultid="43017" />
                    <RANKING order="6" place="6" resultid="41672" />
                    <RANKING order="7" place="-1" resultid="41537" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45396" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42974" />
                    <RANKING order="2" place="2" resultid="43521" />
                    <RANKING order="3" place="-1" resultid="43370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45397" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41697" />
                    <RANKING order="2" place="2" resultid="42102" />
                    <RANKING order="3" place="3" resultid="43131" />
                    <RANKING order="4" place="-1" resultid="41701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45398" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42745" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45399" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41666" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45400" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45401" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45402" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45403" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43822" />
                    <RANKING order="2" place="2" resultid="43946" />
                    <RANKING order="3" place="3" resultid="42050" />
                    <RANKING order="4" place="4" resultid="42821" />
                    <RANKING order="5" place="5" resultid="42779" />
                    <RANKING order="6" place="6" resultid="43893" />
                    <RANKING order="7" place="7" resultid="43919" />
                    <RANKING order="8" place="8" resultid="42012" />
                    <RANKING order="9" place="9" resultid="43085" />
                    <RANKING order="10" place="10" resultid="42989" />
                    <RANKING order="11" place="11" resultid="42974" />
                    <RANKING order="12" place="12" resultid="43943" />
                    <RANKING order="13" place="13" resultid="42868" />
                    <RANKING order="14" place="14" resultid="41877" />
                    <RANKING order="15" place="15" resultid="43307" />
                    <RANKING order="16" place="16" resultid="43135" />
                    <RANKING order="17" place="17" resultid="43365" />
                    <RANKING order="18" place="18" resultid="43675" />
                    <RANKING order="19" place="19" resultid="42677" />
                    <RANKING order="20" place="20" resultid="44008" />
                    <RANKING order="21" place="21" resultid="41910" />
                    <RANKING order="22" place="22" resultid="43346" />
                    <RANKING order="23" place="23" resultid="41983" />
                    <RANKING order="24" place="24" resultid="41810" />
                    <RANKING order="25" place="24" resultid="42476" />
                    <RANKING order="26" place="26" resultid="41697" />
                    <RANKING order="27" place="27" resultid="41967" />
                    <RANKING order="28" place="28" resultid="41900" />
                    <RANKING order="29" place="29" resultid="42191" />
                    <RANKING order="30" place="30" resultid="41739" />
                    <RANKING order="31" place="31" resultid="42181" />
                    <RANKING order="32" place="32" resultid="41719" />
                    <RANKING order="33" place="33" resultid="42019" />
                    <RANKING order="34" place="34" resultid="43463" />
                    <RANKING order="35" place="35" resultid="43888" />
                    <RANKING order="36" place="36" resultid="43076" />
                    <RANKING order="37" place="37" resultid="43532" />
                    <RANKING order="38" place="38" resultid="41834" />
                    <RANKING order="39" place="39" resultid="43521" />
                    <RANKING order="40" place="40" resultid="41751" />
                    <RANKING order="41" place="41" resultid="44854" />
                    <RANKING order="42" place="42" resultid="42001" />
                    <RANKING order="43" place="43" resultid="42102" />
                    <RANKING order="44" place="44" resultid="43980" />
                    <RANKING order="45" place="45" resultid="41860" />
                    <RANKING order="46" place="46" resultid="43409" />
                    <RANKING order="47" place="47" resultid="43131" />
                    <RANKING order="48" place="48" resultid="43017" />
                    <RANKING order="49" place="49" resultid="43696" />
                    <RANKING order="50" place="50" resultid="43839" />
                    <RANKING order="51" place="51" resultid="41666" />
                    <RANKING order="52" place="52" resultid="42745" />
                    <RANKING order="53" place="53" resultid="41672" />
                    <RANKING order="54" place="-1" resultid="43150" />
                    <RANKING order="55" place="-1" resultid="42061" />
                    <RANKING order="56" place="-1" resultid="44003" />
                    <RANKING order="57" place="-1" resultid="41537" />
                    <RANKING order="58" place="-1" resultid="41701" />
                    <RANKING order="59" place="-1" resultid="41830" />
                    <RANKING order="60" place="-1" resultid="42066" />
                    <RANKING order="61" place="-1" resultid="43370" />
                    <RANKING order="62" place="-1" resultid="43468" />
                    <RANKING order="63" place="-1" resultid="43738" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="44975" daytime="16:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="44976" daytime="16:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="44977" daytime="16:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="44978" daytime="16:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="44979" daytime="16:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="44980" daytime="16:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="44981" daytime="16:50" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="44982" daytime="16:55" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2460" daytime="16:55" gender="F" number="21" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45539" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42333" />
                    <RANKING order="2" place="2" resultid="42358" />
                    <RANKING order="3" place="3" resultid="42848" />
                    <RANKING order="4" place="4" resultid="43009" />
                    <RANKING order="5" place="5" resultid="42362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45540" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43081" />
                    <RANKING order="2" place="2" resultid="43775" />
                    <RANKING order="3" place="3" resultid="41544" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45541" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42422" />
                    <RANKING order="2" place="2" resultid="43247" />
                    <RANKING order="3" place="3" resultid="43561" />
                    <RANKING order="4" place="4" resultid="43711" />
                    <RANKING order="5" place="5" resultid="41772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45542" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42733" />
                    <RANKING order="2" place="2" resultid="42509" />
                    <RANKING order="3" place="3" resultid="41549" />
                    <RANKING order="4" place="4" resultid="41623" />
                    <RANKING order="5" place="-1" resultid="43529" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45543" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43872" />
                    <RANKING order="2" place="2" resultid="43242" />
                    <RANKING order="3" place="3" resultid="43198" />
                    <RANKING order="4" place="4" resultid="43626" />
                    <RANKING order="5" place="5" resultid="43232" />
                    <RANKING order="6" place="6" resultid="42760" />
                    <RANKING order="7" place="7" resultid="42842" />
                    <RANKING order="8" place="8" resultid="41816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45544" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42460" />
                    <RANKING order="2" place="2" resultid="43753" />
                    <RANKING order="3" place="3" resultid="44015" />
                    <RANKING order="4" place="4" resultid="42243" />
                    <RANKING order="5" place="-1" resultid="41963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45545" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42073" />
                    <RANKING order="2" place="2" resultid="43976" />
                    <RANKING order="3" place="3" resultid="42969" />
                    <RANKING order="4" place="4" resultid="43878" />
                    <RANKING order="5" place="5" resultid="43748" />
                    <RANKING order="6" place="6" resultid="42407" />
                    <RANKING order="7" place="7" resultid="42825" />
                    <RANKING order="8" place="-1" resultid="43374" />
                    <RANKING order="9" place="-1" resultid="43425" />
                    <RANKING order="10" place="-1" resultid="43867" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45546" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41916" />
                    <RANKING order="2" place="2" resultid="41888" />
                    <RANKING order="3" place="3" resultid="43291" />
                    <RANKING order="4" place="4" resultid="43647" />
                    <RANKING order="5" place="5" resultid="42809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45547" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="43537" />
                    <RANKING order="2" place="-1" resultid="43957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45548" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41820" />
                    <RANKING order="2" place="2" resultid="43228" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45549" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45550" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45551" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45552" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45553" agemax="-1" agemin="-1" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43081" />
                    <RANKING order="2" place="2" resultid="42333" />
                    <RANKING order="3" place="3" resultid="42358" />
                    <RANKING order="4" place="4" resultid="43775" />
                    <RANKING order="5" place="5" resultid="42848" />
                    <RANKING order="6" place="6" resultid="43872" />
                    <RANKING order="7" place="7" resultid="42422" />
                    <RANKING order="8" place="8" resultid="42733" />
                    <RANKING order="9" place="9" resultid="42073" />
                    <RANKING order="10" place="10" resultid="43009" />
                    <RANKING order="11" place="11" resultid="42362" />
                    <RANKING order="12" place="12" resultid="42460" />
                    <RANKING order="13" place="13" resultid="43242" />
                    <RANKING order="14" place="14" resultid="42509" />
                    <RANKING order="15" place="15" resultid="41544" />
                    <RANKING order="16" place="16" resultid="43976" />
                    <RANKING order="17" place="17" resultid="43198" />
                    <RANKING order="18" place="18" resultid="42969" />
                    <RANKING order="19" place="19" resultid="41916" />
                    <RANKING order="20" place="20" resultid="43626" />
                    <RANKING order="21" place="21" resultid="43247" />
                    <RANKING order="22" place="22" resultid="43878" />
                    <RANKING order="23" place="23" resultid="43232" />
                    <RANKING order="24" place="24" resultid="41549" />
                    <RANKING order="25" place="25" resultid="43753" />
                    <RANKING order="26" place="26" resultid="44015" />
                    <RANKING order="27" place="27" resultid="42243" />
                    <RANKING order="28" place="28" resultid="42760" />
                    <RANKING order="29" place="29" resultid="43748" />
                    <RANKING order="30" place="30" resultid="41888" />
                    <RANKING order="31" place="31" resultid="42842" />
                    <RANKING order="32" place="32" resultid="42407" />
                    <RANKING order="33" place="33" resultid="42825" />
                    <RANKING order="34" place="34" resultid="43561" />
                    <RANKING order="35" place="35" resultid="41623" />
                    <RANKING order="36" place="36" resultid="43291" />
                    <RANKING order="37" place="37" resultid="43711" />
                    <RANKING order="38" place="38" resultid="41772" />
                    <RANKING order="39" place="39" resultid="41816" />
                    <RANKING order="40" place="40" resultid="43647" />
                    <RANKING order="41" place="41" resultid="42809" />
                    <RANKING order="42" place="42" resultid="41820" />
                    <RANKING order="43" place="43" resultid="43228" />
                    <RANKING order="44" place="-1" resultid="43374" />
                    <RANKING order="45" place="-1" resultid="43425" />
                    <RANKING order="46" place="-1" resultid="43529" />
                    <RANKING order="47" place="-1" resultid="43537" />
                    <RANKING order="48" place="-1" resultid="43867" />
                    <RANKING order="49" place="-1" resultid="43957" />
                    <RANKING order="50" place="-1" resultid="41963" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45117" daytime="16:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45118" daytime="17:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="45119" daytime="17:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="45120" daytime="17:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="45121" daytime="17:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="45122" daytime="17:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="45123" daytime="17:20" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2445" daytime="17:20" gender="M" number="22" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45374" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43086" />
                    <RANKING order="2" place="-1" resultid="43739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45375" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43931" />
                    <RANKING order="2" place="2" resultid="42780" />
                    <RANKING order="3" place="3" resultid="42013" />
                    <RANKING order="4" place="4" resultid="42711" />
                    <RANKING order="5" place="5" resultid="42434" />
                    <RANKING order="6" place="6" resultid="43786" />
                    <RANKING order="7" place="7" resultid="43151" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45376" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43948" />
                    <RANKING order="2" place="2" resultid="42233" />
                    <RANKING order="3" place="3" resultid="43808" />
                    <RANKING order="4" place="4" resultid="41878" />
                    <RANKING order="5" place="5" resultid="42055" />
                    <RANKING order="6" place="6" resultid="43169" />
                    <RANKING order="7" place="7" resultid="42034" />
                    <RANKING order="8" place="8" resultid="43090" />
                    <RANKING order="9" place="9" resultid="42450" />
                    <RANKING order="10" place="10" resultid="41804" />
                    <RANKING order="11" place="-1" resultid="43145" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45377" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42471" />
                    <RANKING order="2" place="2" resultid="44021" />
                    <RANKING order="3" place="3" resultid="42192" />
                    <RANKING order="4" place="4" resultid="43715" />
                    <RANKING order="5" place="5" resultid="42859" />
                    <RANKING order="6" place="6" resultid="42803" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45378" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41846" />
                    <RANKING order="2" place="2" resultid="42964" />
                    <RANKING order="3" place="3" resultid="41740" />
                    <RANKING order="4" place="4" resultid="41868" />
                    <RANKING order="5" place="5" resultid="42418" />
                    <RANKING order="6" place="6" resultid="43912" />
                    <RANKING order="7" place="7" resultid="43034" />
                    <RANKING order="8" place="8" resultid="43658" />
                    <RANKING order="9" place="-1" resultid="41796" />
                    <RANKING order="10" place="-1" resultid="43443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45379" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43284" />
                    <RANKING order="2" place="2" resultid="42985" />
                    <RANKING order="3" place="3" resultid="41901" />
                    <RANKING order="4" place="4" resultid="42214" />
                    <RANKING order="5" place="5" resultid="42863" />
                    <RANKING order="6" place="6" resultid="43187" />
                    <RANKING order="7" place="7" resultid="43765" />
                    <RANKING order="8" place="8" resultid="41628" />
                    <RANKING order="9" place="9" resultid="43840" />
                    <RANKING order="10" place="10" resultid="43730" />
                    <RANKING order="11" place="11" resultid="42410" />
                    <RANKING order="12" place="12" resultid="43052" />
                    <RANKING order="13" place="-1" resultid="43159" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45380" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43565" />
                    <RANKING order="2" place="2" resultid="43207" />
                    <RANKING order="3" place="3" resultid="42227" />
                    <RANKING order="4" place="4" resultid="42366" />
                    <RANKING order="5" place="5" resultid="41895" />
                    <RANKING order="6" place="6" resultid="42147" />
                    <RANKING order="7" place="7" resultid="43966" />
                    <RANKING order="8" place="8" resultid="42169" />
                    <RANKING order="9" place="-1" resultid="42439" />
                    <RANKING order="10" place="-1" resultid="42756" />
                    <RANKING order="11" place="-1" resultid="42980" />
                    <RANKING order="12" place="-1" resultid="43578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45381" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43216" />
                    <RANKING order="2" place="2" resultid="43884" />
                    <RANKING order="3" place="3" resultid="42129" />
                    <RANKING order="4" place="-1" resultid="43369" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45382" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43266" />
                    <RANKING order="2" place="2" resultid="42496" />
                    <RANKING order="3" place="3" resultid="43393" />
                    <RANKING order="4" place="4" resultid="42154" />
                    <RANKING order="5" place="5" resultid="43154" />
                    <RANKING order="6" place="6" resultid="43496" />
                    <RANKING order="7" place="-1" resultid="41702" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45383" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41872" />
                    <RANKING order="2" place="2" resultid="42415" />
                    <RANKING order="3" place="3" resultid="41679" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45384" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41668" />
                    <RANKING order="2" place="2" resultid="43542" />
                    <RANKING order="3" place="-1" resultid="43582" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45385" agemax="84" agemin="80">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45386" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45387" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45388" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43931" />
                    <RANKING order="2" place="2" resultid="42780" />
                    <RANKING order="3" place="3" resultid="43948" />
                    <RANKING order="4" place="4" resultid="42013" />
                    <RANKING order="5" place="5" resultid="41846" />
                    <RANKING order="6" place="6" resultid="42233" />
                    <RANKING order="7" place="7" resultid="42471" />
                    <RANKING order="8" place="8" resultid="43565" />
                    <RANKING order="9" place="9" resultid="43808" />
                    <RANKING order="10" place="10" resultid="43207" />
                    <RANKING order="11" place="11" resultid="42711" />
                    <RANKING order="12" place="12" resultid="44021" />
                    <RANKING order="13" place="13" resultid="42434" />
                    <RANKING order="14" place="14" resultid="42192" />
                    <RANKING order="15" place="15" resultid="42227" />
                    <RANKING order="16" place="16" resultid="43216" />
                    <RANKING order="17" place="17" resultid="43284" />
                    <RANKING order="18" place="18" resultid="42985" />
                    <RANKING order="19" place="19" resultid="41901" />
                    <RANKING order="20" place="20" resultid="41878" />
                    <RANKING order="21" place="21" resultid="43786" />
                    <RANKING order="22" place="22" resultid="42055" />
                    <RANKING order="23" place="23" resultid="43151" />
                    <RANKING order="24" place="24" resultid="42964" />
                    <RANKING order="25" place="25" resultid="43086" />
                    <RANKING order="26" place="26" resultid="41740" />
                    <RANKING order="27" place="27" resultid="42214" />
                    <RANKING order="28" place="28" resultid="43169" />
                    <RANKING order="29" place="29" resultid="41868" />
                    <RANKING order="30" place="30" resultid="43715" />
                    <RANKING order="31" place="31" resultid="42034" />
                    <RANKING order="32" place="32" resultid="42418" />
                    <RANKING order="33" place="33" resultid="43912" />
                    <RANKING order="34" place="34" resultid="42863" />
                    <RANKING order="35" place="35" resultid="43187" />
                    <RANKING order="36" place="36" resultid="43090" />
                    <RANKING order="37" place="37" resultid="43765" />
                    <RANKING order="38" place="38" resultid="42366" />
                    <RANKING order="39" place="39" resultid="41628" />
                    <RANKING order="40" place="40" resultid="41895" />
                    <RANKING order="41" place="41" resultid="42147" />
                    <RANKING order="42" place="42" resultid="42859" />
                    <RANKING order="43" place="43" resultid="43840" />
                    <RANKING order="44" place="44" resultid="43266" />
                    <RANKING order="45" place="45" resultid="42803" />
                    <RANKING order="46" place="46" resultid="43730" />
                    <RANKING order="47" place="47" resultid="41872" />
                    <RANKING order="48" place="48" resultid="42496" />
                    <RANKING order="49" place="49" resultid="42450" />
                    <RANKING order="50" place="50" resultid="43884" />
                    <RANKING order="51" place="51" resultid="43966" />
                    <RANKING order="52" place="52" resultid="42410" />
                    <RANKING order="53" place="53" resultid="41668" />
                    <RANKING order="54" place="54" resultid="42415" />
                    <RANKING order="55" place="55" resultid="41804" />
                    <RANKING order="56" place="56" resultid="43052" />
                    <RANKING order="57" place="57" resultid="43034" />
                    <RANKING order="58" place="58" resultid="43393" />
                    <RANKING order="59" place="59" resultid="42154" />
                    <RANKING order="60" place="60" resultid="43154" />
                    <RANKING order="61" place="61" resultid="42169" />
                    <RANKING order="62" place="62" resultid="43542" />
                    <RANKING order="63" place="63" resultid="43496" />
                    <RANKING order="64" place="64" resultid="41679" />
                    <RANKING order="65" place="65" resultid="43658" />
                    <RANKING order="66" place="66" resultid="42129" />
                    <RANKING order="67" place="67" resultid="41906" />
                    <RANKING order="68" place="-1" resultid="43159" />
                    <RANKING order="69" place="-1" resultid="42439" />
                    <RANKING order="70" place="-1" resultid="43582" />
                    <RANKING order="71" place="-1" resultid="41702" />
                    <RANKING order="72" place="-1" resultid="41796" />
                    <RANKING order="73" place="-1" resultid="42756" />
                    <RANKING order="74" place="-1" resultid="42980" />
                    <RANKING order="75" place="-1" resultid="43145" />
                    <RANKING order="76" place="-1" resultid="43369" />
                    <RANKING order="77" place="-1" resultid="43443" />
                    <RANKING order="78" place="-1" resultid="43578" />
                    <RANKING order="79" place="-1" resultid="43739" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="44990" daytime="17:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="44991" daytime="17:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="44992" daytime="17:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="44993" daytime="17:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="44994" daytime="17:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="44995" daytime="17:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="44996" daytime="17:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="44997" daytime="17:45" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="44998" daytime="17:45" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="44999" daytime="17:50" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2021-07-11" daytime="09:30" endtime="12:19" name="3ª Jornada-1ª sessão" number="5">
          <EVENTS>
            <EVENT eventid="2263" daytime="09:30" gender="M" number="23" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45359" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42371" />
                    <RANKING order="2" place="2" resultid="42815" />
                    <RANKING order="3" place="3" resultid="43601" />
                    <RANKING order="4" place="4" resultid="43705" />
                    <RANKING order="5" place="5" resultid="41735" />
                    <RANKING order="6" place="6" resultid="43486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45360" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43826" />
                    <RANKING order="2" place="2" resultid="43309" />
                    <RANKING order="3" place="3" resultid="43136" />
                    <RANKING order="4" place="-1" resultid="43861" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45361" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43474" />
                    <RANKING order="2" place="2" resultid="42006" />
                    <RANKING order="3" place="3" resultid="44009" />
                    <RANKING order="4" place="4" resultid="43077" />
                    <RANKING order="5" place="5" resultid="42062" />
                    <RANKING order="6" place="6" resultid="42035" />
                    <RANKING order="7" place="7" resultid="43091" />
                    <RANKING order="8" place="8" resultid="43410" />
                    <RANKING order="9" place="-1" resultid="41831" />
                    <RANKING order="10" place="-1" resultid="43170" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45362" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42089" />
                    <RANKING order="2" place="2" resultid="42764" />
                    <RANKING order="3" place="3" resultid="42067" />
                    <RANKING order="4" place="4" resultid="42424" />
                    <RANKING order="5" place="5" resultid="43697" />
                    <RANKING order="6" place="-1" resultid="43404" />
                    <RANKING order="7" place="-1" resultid="41958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45363" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43176" />
                    <RANKING order="2" place="2" resultid="41968" />
                    <RANKING order="3" place="3" resultid="43599" />
                    <RANKING order="4" place="4" resultid="42095" />
                    <RANKING order="5" place="5" resultid="42957" />
                    <RANKING order="6" place="6" resultid="43691" />
                    <RANKING order="7" place="-1" resultid="42428" />
                    <RANKING order="8" place="-1" resultid="43996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45364" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41902" />
                    <RANKING order="2" place="2" resultid="43764" />
                    <RANKING order="3" place="3" resultid="43835" />
                    <RANKING order="4" place="4" resultid="43352" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45365" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43613" />
                    <RANKING order="2" place="2" resultid="43551" />
                    <RANKING order="3" place="3" resultid="43193" />
                    <RANKING order="4" place="4" resultid="41861" />
                    <RANKING order="5" place="5" resultid="43072" />
                    <RANKING order="6" place="6" resultid="42167" />
                    <RANKING order="7" place="-1" resultid="43208" />
                    <RANKING order="8" place="-1" resultid="43555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45366" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41687" />
                    <RANKING order="2" place="2" resultid="43217" />
                    <RANKING order="3" place="3" resultid="43522" />
                    <RANKING order="4" place="4" resultid="43883" />
                    <RANKING order="5" place="5" resultid="43491" />
                    <RANKING order="6" place="6" resultid="43453" />
                    <RANKING order="7" place="-1" resultid="43371" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45367" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43132" />
                    <RANKING order="2" place="2" resultid="42752" />
                    <RANKING order="3" place="3" resultid="42495" />
                    <RANKING order="4" place="4" resultid="41765" />
                    <RANKING order="5" place="5" resultid="43028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45368" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41662" />
                    <RANKING order="2" place="2" resultid="41678" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45369" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45370" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45371" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45372" agemax="94" agemin="90">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="41852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45373" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43826" />
                    <RANKING order="2" place="2" resultid="43613" />
                    <RANKING order="3" place="3" resultid="43474" />
                    <RANKING order="4" place="4" resultid="43176" />
                    <RANKING order="5" place="5" resultid="42089" />
                    <RANKING order="6" place="6" resultid="42371" />
                    <RANKING order="7" place="7" resultid="42764" />
                    <RANKING order="8" place="8" resultid="42815" />
                    <RANKING order="9" place="9" resultid="42006" />
                    <RANKING order="10" place="10" resultid="43309" />
                    <RANKING order="11" place="11" resultid="41687" />
                    <RANKING order="12" place="12" resultid="43601" />
                    <RANKING order="13" place="13" resultid="41968" />
                    <RANKING order="14" place="14" resultid="44009" />
                    <RANKING order="15" place="15" resultid="43705" />
                    <RANKING order="16" place="16" resultid="43599" />
                    <RANKING order="17" place="17" resultid="42095" />
                    <RANKING order="18" place="18" resultid="42957" />
                    <RANKING order="19" place="19" resultid="41735" />
                    <RANKING order="20" place="20" resultid="43136" />
                    <RANKING order="21" place="21" resultid="43691" />
                    <RANKING order="22" place="22" resultid="43217" />
                    <RANKING order="23" place="23" resultid="41902" />
                    <RANKING order="24" place="24" resultid="42067" />
                    <RANKING order="25" place="25" resultid="43522" />
                    <RANKING order="26" place="26" resultid="41662" />
                    <RANKING order="27" place="27" resultid="43077" />
                    <RANKING order="28" place="28" resultid="42424" />
                    <RANKING order="29" place="29" resultid="43551" />
                    <RANKING order="30" place="30" resultid="42062" />
                    <RANKING order="31" place="31" resultid="42035" />
                    <RANKING order="32" place="32" resultid="43697" />
                    <RANKING order="33" place="33" resultid="43193" />
                    <RANKING order="34" place="34" resultid="43091" />
                    <RANKING order="35" place="35" resultid="43764" />
                    <RANKING order="36" place="36" resultid="43132" />
                    <RANKING order="37" place="37" resultid="41861" />
                    <RANKING order="38" place="38" resultid="43072" />
                    <RANKING order="39" place="39" resultid="42752" />
                    <RANKING order="40" place="40" resultid="43835" />
                    <RANKING order="41" place="41" resultid="43883" />
                    <RANKING order="42" place="42" resultid="43491" />
                    <RANKING order="43" place="43" resultid="42495" />
                    <RANKING order="44" place="44" resultid="43352" />
                    <RANKING order="45" place="45" resultid="41765" />
                    <RANKING order="46" place="46" resultid="43028" />
                    <RANKING order="47" place="47" resultid="43486" />
                    <RANKING order="48" place="48" resultid="42167" />
                    <RANKING order="49" place="49" resultid="41655" />
                    <RANKING order="50" place="50" resultid="43410" />
                    <RANKING order="51" place="51" resultid="43453" />
                    <RANKING order="52" place="52" resultid="41678" />
                    <RANKING order="53" place="-1" resultid="41831" />
                    <RANKING order="54" place="-1" resultid="41852" />
                    <RANKING order="55" place="-1" resultid="42428" />
                    <RANKING order="56" place="-1" resultid="43170" />
                    <RANKING order="57" place="-1" resultid="43208" />
                    <RANKING order="58" place="-1" resultid="43371" />
                    <RANKING order="59" place="-1" resultid="43404" />
                    <RANKING order="60" place="-1" resultid="43555" />
                    <RANKING order="61" place="-1" resultid="43861" />
                    <RANKING order="62" place="-1" resultid="41958" />
                    <RANKING order="63" place="-1" resultid="43996" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45124" daytime="09:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45125" daytime="09:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="45126" daytime="09:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="45127" daytime="10:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="45128" daytime="10:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="45129" daytime="10:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="45130" daytime="10:25" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="45131" daytime="10:30" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2492" daytime="10:40" gender="F" number="24" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45524" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42996" />
                    <RANKING order="2" place="2" resultid="42455" />
                    <RANKING order="3" place="3" resultid="42465" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45525" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43663" />
                    <RANKING order="2" place="2" resultid="41543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45526" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41995" />
                    <RANKING order="2" place="2" resultid="42238" />
                    <RANKING order="3" place="3" resultid="43312" />
                    <RANKING order="4" place="4" resultid="43248" />
                    <RANKING order="5" place="5" resultid="41773" />
                    <RANKING order="6" place="-1" resultid="42445" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45527" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43066" />
                    <RANKING order="2" place="2" resultid="42698" />
                    <RANKING order="3" place="3" resultid="43907" />
                    <RANKING order="4" place="4" resultid="42508" />
                    <RANKING order="5" place="5" resultid="43272" />
                    <RANKING order="6" place="6" resultid="43400" />
                    <RANKING order="7" place="7" resultid="43337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45528" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42122" />
                    <RANKING order="2" place="2" resultid="43500" />
                    <RANKING order="3" place="3" resultid="42031" />
                    <RANKING order="4" place="4" resultid="41946" />
                    <RANKING order="5" place="5" resultid="43354" />
                    <RANKING order="6" place="-1" resultid="43199" />
                    <RANKING order="7" place="-1" resultid="43769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45529" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42047" />
                    <RANKING order="2" place="2" resultid="43222" />
                    <RANKING order="3" place="3" resultid="43433" />
                    <RANKING order="4" place="4" resultid="42176" />
                    <RANKING order="5" place="5" resultid="43681" />
                    <RANKING order="6" place="6" resultid="41938" />
                    <RANKING order="7" place="7" resultid="44016" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45530" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43975" />
                    <RANKING order="2" place="2" resultid="42970" />
                    <RANKING order="3" place="3" resultid="41922" />
                    <RANKING order="4" place="4" resultid="43877" />
                    <RANKING order="5" place="5" resultid="42208" />
                    <RANKING order="6" place="6" resultid="43866" />
                    <RANKING order="7" place="7" resultid="43126" />
                    <RANKING order="8" place="8" resultid="42692" />
                    <RANKING order="9" place="-1" resultid="43426" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45531" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43852" />
                    <RANKING order="2" place="2" resultid="41747" />
                    <RANKING order="3" place="3" resultid="43292" />
                    <RANKING order="4" place="-1" resultid="43572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45532" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="45533" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="45534" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45535" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45536" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45537" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45538" agemax="-1" agemin="-1" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42996" />
                    <RANKING order="2" place="2" resultid="42455" />
                    <RANKING order="3" place="3" resultid="41995" />
                    <RANKING order="4" place="4" resultid="42122" />
                    <RANKING order="5" place="5" resultid="43663" />
                    <RANKING order="6" place="6" resultid="42047" />
                    <RANKING order="7" place="7" resultid="43066" />
                    <RANKING order="8" place="8" resultid="43222" />
                    <RANKING order="9" place="9" resultid="42698" />
                    <RANKING order="10" place="10" resultid="43907" />
                    <RANKING order="11" place="11" resultid="43500" />
                    <RANKING order="12" place="12" resultid="42508" />
                    <RANKING order="13" place="13" resultid="41543" />
                    <RANKING order="14" place="14" resultid="42465" />
                    <RANKING order="15" place="15" resultid="43272" />
                    <RANKING order="16" place="16" resultid="43433" />
                    <RANKING order="17" place="17" resultid="43975" />
                    <RANKING order="18" place="18" resultid="42970" />
                    <RANKING order="19" place="19" resultid="41922" />
                    <RANKING order="20" place="20" resultid="43877" />
                    <RANKING order="21" place="21" resultid="43400" />
                    <RANKING order="22" place="22" resultid="42208" />
                    <RANKING order="23" place="23" resultid="42031" />
                    <RANKING order="24" place="24" resultid="42176" />
                    <RANKING order="25" place="25" resultid="43866" />
                    <RANKING order="26" place="26" resultid="43852" />
                    <RANKING order="27" place="27" resultid="42238" />
                    <RANKING order="28" place="28" resultid="43681" />
                    <RANKING order="29" place="29" resultid="41938" />
                    <RANKING order="30" place="30" resultid="43126" />
                    <RANKING order="31" place="31" resultid="41946" />
                    <RANKING order="32" place="32" resultid="42692" />
                    <RANKING order="33" place="33" resultid="43312" />
                    <RANKING order="34" place="34" resultid="44016" />
                    <RANKING order="35" place="35" resultid="41747" />
                    <RANKING order="36" place="36" resultid="43248" />
                    <RANKING order="37" place="37" resultid="41773" />
                    <RANKING order="38" place="38" resultid="43337" />
                    <RANKING order="39" place="39" resultid="43292" />
                    <RANKING order="40" place="40" resultid="43354" />
                    <RANKING order="41" place="-1" resultid="42445" />
                    <RANKING order="42" place="-1" resultid="43199" />
                    <RANKING order="43" place="-1" resultid="43426" />
                    <RANKING order="44" place="-1" resultid="43572" />
                    <RANKING order="45" place="-1" resultid="43769" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45008" daytime="10:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45009" daytime="10:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="45010" daytime="11:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="45011" daytime="11:05" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="45012" daytime="11:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="45013" daytime="11:25" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2293" daytime="11:30" gender="M" number="25" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45344" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41825" />
                    <RANKING order="2" place="2" resultid="42704" />
                    <RANKING order="3" place="3" resultid="42836" />
                    <RANKING order="4" place="4" resultid="43602" />
                    <RANKING order="5" place="5" resultid="42798" />
                    <RANKING order="6" place="6" resultid="42376" />
                    <RANKING order="7" place="7" resultid="43605" />
                    <RANKING order="8" place="8" resultid="42678" />
                    <RANKING order="9" place="9" resultid="43341" />
                    <RANKING order="10" place="-1" resultid="42342" />
                    <RANKING order="11" place="-1" resultid="42789" />
                    <RANKING order="12" place="-1" resultid="43201" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45345" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42106" />
                    <RANKING order="2" place="2" resultid="43164" />
                    <RANKING order="3" place="3" resultid="41952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45346" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43947" />
                    <RANKING order="2" place="2" resultid="43920" />
                    <RANKING order="3" place="3" resultid="41648" />
                    <RANKING order="4" place="3" resultid="44855" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45347" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43469" />
                    <RANKING order="2" place="2" resultid="43366" />
                    <RANKING order="3" place="3" resultid="42068" />
                    <RANKING order="4" place="4" resultid="43796" />
                    <RANKING order="5" place="5" resultid="41839" />
                    <RANKING order="6" place="6" resultid="42248" />
                    <RANKING order="7" place="7" resultid="44004" />
                    <RANKING order="8" place="8" resultid="42804" />
                    <RANKING order="9" place="9" resultid="43981" />
                    <RANKING order="10" place="-1" resultid="41728" />
                    <RANKING order="11" place="-1" resultid="43735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45348" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43588" />
                    <RANKING order="2" place="2" resultid="42480" />
                    <RANKING order="3" place="3" resultid="43379" />
                    <RANKING order="4" place="4" resultid="42830" />
                    <RANKING order="5" place="5" resultid="43033" />
                    <RANKING order="6" place="6" resultid="43657" />
                    <RANKING order="7" place="-1" resultid="41619" />
                    <RANKING order="8" place="-1" resultid="43998" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45349" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42220" />
                    <RANKING order="2" place="2" resultid="43387" />
                    <RANKING order="3" place="3" resultid="42490" />
                    <RANKING order="4" place="4" resultid="41635" />
                    <RANKING order="5" place="5" resultid="43889" />
                    <RANKING order="6" place="6" resultid="42722" />
                    <RANKING order="7" place="7" resultid="43506" />
                    <RANKING order="8" place="-1" resultid="42112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45350" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42226" />
                    <RANKING order="2" place="2" resultid="43347" />
                    <RANKING order="3" place="3" resultid="43566" />
                    <RANKING order="4" place="4" resultid="43059" />
                    <RANKING order="5" place="5" resultid="43926" />
                    <RANKING order="6" place="6" resultid="41896" />
                    <RANKING order="7" place="7" resultid="43552" />
                    <RANKING order="8" place="8" resultid="42680" />
                    <RANKING order="9" place="9" resultid="43965" />
                    <RANKING order="10" place="10" resultid="42168" />
                    <RANKING order="11" place="-1" resultid="43510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45351" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43516" />
                    <RANKING order="2" place="2" resultid="42117" />
                    <RANKING order="3" place="3" resultid="42040" />
                    <RANKING order="4" place="4" resultid="42128" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45352" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43267" />
                    <RANKING order="2" place="2" resultid="43394" />
                    <RANKING order="3" place="3" resultid="43029" />
                    <RANKING order="4" place="4" resultid="42153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45353" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41873" />
                    <RANKING order="2" place="2" resultid="43360" />
                    <RANKING order="3" place="3" resultid="42746" />
                    <RANKING order="4" place="-1" resultid="41713" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45354" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41667" />
                    <RANKING order="2" place="2" resultid="43543" />
                    <RANKING order="3" place="3" resultid="43583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45355" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45356" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45357" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45358" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41825" />
                    <RANKING order="2" place="2" resultid="42704" />
                    <RANKING order="3" place="3" resultid="42106" />
                    <RANKING order="4" place="4" resultid="42220" />
                    <RANKING order="5" place="5" resultid="43947" />
                    <RANKING order="6" place="6" resultid="43920" />
                    <RANKING order="7" place="7" resultid="43588" />
                    <RANKING order="8" place="8" resultid="42836" />
                    <RANKING order="9" place="8" resultid="43387" />
                    <RANKING order="10" place="10" resultid="43602" />
                    <RANKING order="11" place="11" resultid="43469" />
                    <RANKING order="12" place="12" resultid="42798" />
                    <RANKING order="13" place="13" resultid="42376" />
                    <RANKING order="14" place="14" resultid="42490" />
                    <RANKING order="15" place="15" resultid="41635" />
                    <RANKING order="16" place="16" resultid="42480" />
                    <RANKING order="17" place="17" resultid="43605" />
                    <RANKING order="18" place="18" resultid="42226" />
                    <RANKING order="19" place="19" resultid="42678" />
                    <RANKING order="20" place="20" resultid="43347" />
                    <RANKING order="21" place="21" resultid="43341" />
                    <RANKING order="22" place="22" resultid="43366" />
                    <RANKING order="23" place="23" resultid="43889" />
                    <RANKING order="24" place="24" resultid="42068" />
                    <RANKING order="25" place="25" resultid="43796" />
                    <RANKING order="26" place="26" resultid="41839" />
                    <RANKING order="27" place="27" resultid="43566" />
                    <RANKING order="28" place="28" resultid="43379" />
                    <RANKING order="29" place="29" resultid="43164" />
                    <RANKING order="30" place="30" resultid="43516" />
                    <RANKING order="31" place="31" resultid="42722" />
                    <RANKING order="32" place="32" resultid="42248" />
                    <RANKING order="33" place="33" resultid="43506" />
                    <RANKING order="34" place="34" resultid="43059" />
                    <RANKING order="35" place="35" resultid="43926" />
                    <RANKING order="36" place="36" resultid="42117" />
                    <RANKING order="37" place="37" resultid="41648" />
                    <RANKING order="38" place="37" resultid="44855" />
                    <RANKING order="39" place="39" resultid="41952" />
                    <RANKING order="40" place="40" resultid="41896" />
                    <RANKING order="41" place="41" resultid="43552" />
                    <RANKING order="42" place="42" resultid="42830" />
                    <RANKING order="43" place="43" resultid="44004" />
                    <RANKING order="44" place="44" resultid="42804" />
                    <RANKING order="45" place="45" resultid="42040" />
                    <RANKING order="46" place="46" resultid="43267" />
                    <RANKING order="47" place="47" resultid="43033" />
                    <RANKING order="48" place="48" resultid="41873" />
                    <RANKING order="49" place="49" resultid="43981" />
                    <RANKING order="50" place="50" resultid="43394" />
                    <RANKING order="51" place="51" resultid="42680" />
                    <RANKING order="52" place="52" resultid="43029" />
                    <RANKING order="53" place="53" resultid="43965" />
                    <RANKING order="54" place="54" resultid="41667" />
                    <RANKING order="55" place="55" resultid="43360" />
                    <RANKING order="56" place="56" resultid="42746" />
                    <RANKING order="57" place="57" resultid="43657" />
                    <RANKING order="58" place="58" resultid="43543" />
                    <RANKING order="59" place="59" resultid="43583" />
                    <RANKING order="60" place="60" resultid="42153" />
                    <RANKING order="61" place="61" resultid="42168" />
                    <RANKING order="62" place="62" resultid="42128" />
                    <RANKING order="63" place="-1" resultid="41619" />
                    <RANKING order="64" place="-1" resultid="41713" />
                    <RANKING order="65" place="-1" resultid="41728" />
                    <RANKING order="66" place="-1" resultid="42112" />
                    <RANKING order="67" place="-1" resultid="42342" />
                    <RANKING order="68" place="-1" resultid="42789" />
                    <RANKING order="69" place="-1" resultid="43201" />
                    <RANKING order="70" place="-1" resultid="43510" />
                    <RANKING order="71" place="-1" resultid="43735" />
                    <RANKING order="72" place="-1" resultid="43998" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45014" daytime="11:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45015" daytime="11:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="45016" daytime="11:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="45017" daytime="11:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="45018" daytime="11:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="45019" daytime="11:45" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="45020" daytime="11:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="45021" daytime="11:50" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="45022" daytime="11:50" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2522" daytime="11:55" gender="F" number="26" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45509" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42785" />
                    <RANKING order="2" place="2" resultid="42739" />
                    <RANKING order="3" place="3" resultid="42159" />
                    <RANKING order="4" place="4" resultid="42345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45510" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43970" />
                    <RANKING order="2" place="2" resultid="43638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45511" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41996" />
                    <RANKING order="2" place="2" resultid="43414" />
                    <RANKING order="3" place="3" resultid="43780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45512" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43846" />
                    <RANKING order="2" place="2" resultid="43041" />
                    <RANKING order="3" place="3" resultid="43273" />
                    <RANKING order="4" place="4" resultid="43908" />
                    <RANKING order="5" place="5" resultid="42852" />
                    <RANKING order="6" place="6" resultid="42726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45513" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42123" />
                    <RANKING order="2" place="2" resultid="43829" />
                    <RANKING order="3" place="3" resultid="41990" />
                    <RANKING order="4" place="4" resultid="43253" />
                    <RANKING order="5" place="5" resultid="42716" />
                    <RANKING order="6" place="6" resultid="43458" />
                    <RANKING order="7" place="-1" resultid="43595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45514" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43303" />
                    <RANKING order="2" place="2" resultid="43431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45515" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42141" />
                    <RANKING order="2" place="2" resultid="43438" />
                    <RANKING order="3" place="3" resultid="42072" />
                    <RANKING order="4" place="4" resultid="42209" />
                    <RANKING order="5" place="5" resultid="43939" />
                    <RANKING order="6" place="6" resultid="43237" />
                    <RANKING order="7" place="7" resultid="43480" />
                    <RANKING order="8" place="-1" resultid="43427" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45516" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41704" />
                    <RANKING order="2" place="2" resultid="42810" />
                    <RANKING order="3" place="3" resultid="41889" />
                    <RANKING order="4" place="4" resultid="43140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45517" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41883" />
                    <RANKING order="2" place="2" resultid="43956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45518" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41821" />
                    <RANKING order="2" place="-1" resultid="41707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45519" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45520" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45521" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45522" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45523" agemax="-1" agemin="-1" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42785" />
                    <RANKING order="2" place="2" resultid="42739" />
                    <RANKING order="3" place="3" resultid="43970" />
                    <RANKING order="4" place="4" resultid="43846" />
                    <RANKING order="5" place="5" resultid="42123" />
                    <RANKING order="6" place="6" resultid="41996" />
                    <RANKING order="7" place="7" resultid="42159" />
                    <RANKING order="8" place="8" resultid="42345" />
                    <RANKING order="9" place="9" resultid="43414" />
                    <RANKING order="10" place="10" resultid="43041" />
                    <RANKING order="11" place="11" resultid="43303" />
                    <RANKING order="12" place="12" resultid="43638" />
                    <RANKING order="13" place="13" resultid="42141" />
                    <RANKING order="14" place="14" resultid="43829" />
                    <RANKING order="15" place="15" resultid="43780" />
                    <RANKING order="16" place="16" resultid="43438" />
                    <RANKING order="17" place="17" resultid="42072" />
                    <RANKING order="18" place="18" resultid="43273" />
                    <RANKING order="19" place="19" resultid="41990" />
                    <RANKING order="20" place="20" resultid="43908" />
                    <RANKING order="21" place="21" resultid="41704" />
                    <RANKING order="22" place="22" resultid="42852" />
                    <RANKING order="23" place="23" resultid="43431" />
                    <RANKING order="24" place="24" resultid="43253" />
                    <RANKING order="25" place="25" resultid="42716" />
                    <RANKING order="26" place="26" resultid="42726" />
                    <RANKING order="27" place="27" resultid="42209" />
                    <RANKING order="28" place="28" resultid="43939" />
                    <RANKING order="29" place="29" resultid="43458" />
                    <RANKING order="30" place="30" resultid="43237" />
                    <RANKING order="31" place="31" resultid="41883" />
                    <RANKING order="32" place="32" resultid="42810" />
                    <RANKING order="33" place="33" resultid="41889" />
                    <RANKING order="34" place="34" resultid="43480" />
                    <RANKING order="35" place="35" resultid="43140" />
                    <RANKING order="36" place="36" resultid="41821" />
                    <RANKING order="37" place="37" resultid="43956" />
                    <RANKING order="38" place="-1" resultid="41707" />
                    <RANKING order="39" place="-1" resultid="43427" />
                    <RANKING order="40" place="-1" resultid="43595" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45023" daytime="11:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45024" daytime="11:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="45025" daytime="12:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="45026" daytime="12:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="45027" daytime="12:05" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2567" daytime="12:05" gender="M" number="27" order="5" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45329" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41799" />
                    <RANKING order="2" place="-1" resultid="42327" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45330" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45331" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43823" />
                    <RANKING order="2" place="2" resultid="42007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45332" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42990" />
                    <RANKING order="2" place="2" resultid="42090" />
                    <RANKING order="3" place="3" resultid="41911" />
                    <RANKING order="4" place="4" resultid="41752" />
                    <RANKING order="5" place="-1" resultid="43464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45333" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41792" />
                    <RANKING order="2" place="2" resultid="42096" />
                    <RANKING order="3" place="3" resultid="43421" />
                    <RANKING order="4" place="4" resultid="43449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45334" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42477" />
                    <RANKING order="2" place="2" resultid="42182" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45335" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43344" />
                    <RANKING order="2" place="-1" resultid="42002" />
                    <RANKING order="3" place="-1" resultid="41673" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45336" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42975" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45337" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43022" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45338" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="45339" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45340" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45341" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45342" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45343" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41799" />
                    <RANKING order="2" place="2" resultid="43823" />
                    <RANKING order="3" place="3" resultid="42975" />
                    <RANKING order="4" place="4" resultid="42990" />
                    <RANKING order="5" place="5" resultid="41792" />
                    <RANKING order="6" place="6" resultid="42007" />
                    <RANKING order="7" place="7" resultid="43137" />
                    <RANKING order="8" place="8" resultid="42090" />
                    <RANKING order="9" place="9" resultid="42477" />
                    <RANKING order="10" place="10" resultid="41911" />
                    <RANKING order="11" place="11" resultid="42182" />
                    <RANKING order="12" place="12" resultid="42096" />
                    <RANKING order="13" place="13" resultid="43344" />
                    <RANKING order="14" place="14" resultid="43421" />
                    <RANKING order="15" place="15" resultid="41752" />
                    <RANKING order="16" place="16" resultid="43449" />
                    <RANKING order="17" place="17" resultid="43022" />
                    <RANKING order="18" place="-1" resultid="42002" />
                    <RANKING order="19" place="-1" resultid="41673" />
                    <RANKING order="20" place="-1" resultid="43464" />
                    <RANKING order="21" place="-1" resultid="42327" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45028" daytime="12:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45029" daytime="12:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="45030" daytime="12:20" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2667" daytime="12:25" gender="F" number="28" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45494" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="44031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45495" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45496" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="43249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45497" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="45498" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43871" />
                    <RANKING order="2" place="2" resultid="43254" />
                    <RANKING order="3" place="3" resultid="43355" />
                    <RANKING order="4" place="-1" resultid="43770" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45499" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="45500" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45501" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="45502" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="45503" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="45504" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45505" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45506" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45507" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45508" agemax="-1" agemin="-1" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41725" />
                    <RANKING order="2" place="2" resultid="44031" />
                    <RANKING order="3" place="3" resultid="43871" />
                    <RANKING order="4" place="4" resultid="43254" />
                    <RANKING order="5" place="5" resultid="42136" />
                    <RANKING order="6" place="6" resultid="43355" />
                    <RANKING order="7" place="-1" resultid="43249" />
                    <RANKING order="8" place="-1" resultid="43770" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45031" daytime="12:25" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2021-07-11" daytime="15:30" endtime="17:15" name="3ª Jornada-2ª sessão" number="6">
          <EVENTS>
            <EVENT eventid="2652" daytime="15:30" gender="M" number="29" order="1" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45314" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42328" />
                    <RANKING order="2" place="2" resultid="42822" />
                    <RANKING order="3" place="3" resultid="43202" />
                    <RANKING order="4" place="4" resultid="43936" />
                    <RANKING order="5" place="5" resultid="42837" />
                    <RANKING order="6" place="6" resultid="42372" />
                    <RANKING order="7" place="7" resultid="42670" />
                    <RANKING order="8" place="8" resultid="42799" />
                    <RANKING order="9" place="9" resultid="42816" />
                    <RANKING order="10" place="10" resultid="43606" />
                    <RANKING order="11" place="11" resultid="42377" />
                    <RANKING order="12" place="12" resultid="42687" />
                    <RANKING order="13" place="13" resultid="42869" />
                    <RANKING order="14" place="14" resultid="43706" />
                    <RANKING order="15" place="-1" resultid="41826" />
                    <RANKING order="16" place="-1" resultid="42343" />
                    <RANKING order="17" place="-1" resultid="43002" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45315" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42107" />
                    <RANKING order="2" place="2" resultid="43745" />
                    <RANKING order="3" place="3" resultid="43894" />
                    <RANKING order="4" place="4" resultid="42435" />
                    <RANKING order="5" place="5" resultid="43676" />
                    <RANKING order="6" place="6" resultid="43655" />
                    <RANKING order="7" place="7" resultid="43787" />
                    <RANKING order="8" place="8" resultid="41953" />
                    <RANKING order="9" place="9" resultid="43165" />
                    <RANKING order="10" place="-1" resultid="41532" />
                    <RANKING order="11" place="-1" resultid="42026" />
                    <RANKING order="12" place="-1" resultid="42348" />
                    <RANKING order="13" place="-1" resultid="43270" />
                    <RANKING order="14" place="-1" resultid="43862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45316" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42773" />
                    <RANKING order="2" place="2" resultid="43475" />
                    <RANKING order="3" place="3" resultid="43004" />
                    <RANKING order="4" place="4" resultid="42486" />
                    <RANKING order="5" place="5" resultid="43921" />
                    <RANKING order="6" place="6" resultid="41879" />
                    <RANKING order="7" place="7" resultid="43814" />
                    <RANKING order="8" place="8" resultid="43701" />
                    <RANKING order="9" place="9" resultid="44010" />
                    <RANKING order="10" place="10" resultid="42056" />
                    <RANKING order="11" place="11" resultid="41649" />
                    <RANKING order="12" place="12" resultid="41805" />
                    <RANKING order="13" place="-1" resultid="43146" />
                    <RANKING order="14" place="-1" resultid="43171" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45317" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43470" />
                    <RANKING order="2" place="2" resultid="42091" />
                    <RANKING order="3" place="3" resultid="43367" />
                    <RANKING order="4" place="4" resultid="42729" />
                    <RANKING order="5" place="5" resultid="42472" />
                    <RANKING order="6" place="6" resultid="43797" />
                    <RANKING order="7" place="7" resultid="41840" />
                    <RANKING order="8" place="8" resultid="42249" />
                    <RANKING order="9" place="9" resultid="44022" />
                    <RANKING order="10" place="10" resultid="43688" />
                    <RANKING order="11" place="11" resultid="43982" />
                    <RANKING order="12" place="12" resultid="43734" />
                    <RANKING order="13" place="13" resultid="41753" />
                    <RANKING order="14" place="14" resultid="42805" />
                    <RANKING order="15" place="15" resultid="44005" />
                    <RANKING order="16" place="16" resultid="43716" />
                    <RANKING order="17" place="-1" resultid="41925" />
                    <RANKING order="18" place="-1" resultid="41729" />
                    <RANKING order="19" place="-1" resultid="42336" />
                    <RANKING order="20" place="-1" resultid="42425" />
                    <RANKING order="21" place="-1" resultid="41521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45318" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43177" />
                    <RANKING order="2" place="2" resultid="42481" />
                    <RANKING order="3" place="3" resultid="42965" />
                    <RANKING order="4" place="4" resultid="43380" />
                    <RANKING order="5" place="5" resultid="42958" />
                    <RANKING order="6" place="6" resultid="43992" />
                    <RANKING order="7" place="7" resultid="42831" />
                    <RANKING order="8" place="8" resultid="43035" />
                    <RANKING order="9" place="9" resultid="43913" />
                    <RANKING order="10" place="10" resultid="43725" />
                    <RANKING order="11" place="-1" resultid="43629" />
                    <RANKING order="12" place="-1" resultid="43856" />
                    <RANKING order="13" place="-1" resultid="43999" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45319" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42221" />
                    <RANKING order="2" place="2" resultid="43388" />
                    <RANKING order="3" place="3" resultid="42491" />
                    <RANKING order="4" place="4" resultid="41636" />
                    <RANKING order="5" place="5" resultid="43260" />
                    <RANKING order="6" place="6" resultid="43890" />
                    <RANKING order="7" place="7" resultid="42215" />
                    <RANKING order="8" place="8" resultid="43006" />
                    <RANKING order="9" place="9" resultid="43286" />
                    <RANKING order="10" place="10" resultid="42723" />
                    <RANKING order="11" place="11" resultid="44026" />
                    <RANKING order="12" place="12" resultid="43593" />
                    <RANKING order="13" place="13" resultid="43671" />
                    <RANKING order="14" place="14" resultid="43731" />
                    <RANKING order="15" place="15" resultid="42672" />
                    <RANKING order="16" place="16" resultid="43160" />
                    <RANKING order="17" place="-1" resultid="42792" />
                    <RANKING order="18" place="-1" resultid="43383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45320" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41720" />
                    <RANKING order="2" place="2" resultid="43927" />
                    <RANKING order="3" place="3" resultid="43553" />
                    <RANKING order="4" place="4" resultid="43060" />
                    <RANKING order="5" place="5" resultid="42367" />
                    <RANKING order="6" place="6" resultid="42148" />
                    <RANKING order="7" place="7" resultid="41862" />
                    <RANKING order="8" place="8" resultid="42681" />
                    <RANKING order="9" place="9" resultid="43621" />
                    <RANKING order="10" place="10" resultid="43073" />
                    <RANKING order="11" place="-1" resultid="43567" />
                    <RANKING order="12" place="-1" resultid="43511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45321" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41688" />
                    <RANKING order="2" place="2" resultid="43517" />
                    <RANKING order="3" place="3" resultid="42118" />
                    <RANKING order="4" place="4" resultid="42041" />
                    <RANKING order="5" place="5" resultid="42130" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45322" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41766" />
                    <RANKING order="2" place="2" resultid="43395" />
                    <RANKING order="3" place="3" resultid="42753" />
                    <RANKING order="4" place="4" resultid="43023" />
                    <RANKING order="5" place="5" resultid="43497" />
                    <RANKING order="6" place="6" resultid="43155" />
                    <RANKING order="7" place="-1" resultid="42497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45323" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41682" />
                    <RANKING order="2" place="2" resultid="41874" />
                    <RANKING order="3" place="3" resultid="43361" />
                    <RANKING order="4" place="4" resultid="41680" />
                    <RANKING order="5" place="5" resultid="42404" />
                    <RANKING order="6" place="-1" resultid="41714" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45324" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41656" />
                    <RANKING order="2" place="2" resultid="43584" />
                    <RANKING order="3" place="3" resultid="43544" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45325" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45326" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45327" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45328" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42107" />
                    <RANKING order="2" place="2" resultid="42773" />
                    <RANKING order="3" place="3" resultid="42328" />
                    <RANKING order="4" place="4" resultid="42822" />
                    <RANKING order="5" place="5" resultid="43745" />
                    <RANKING order="6" place="6" resultid="43202" />
                    <RANKING order="7" place="7" resultid="43475" />
                    <RANKING order="8" place="8" resultid="43936" />
                    <RANKING order="9" place="9" resultid="42837" />
                    <RANKING order="10" place="10" resultid="42372" />
                    <RANKING order="11" place="11" resultid="43894" />
                    <RANKING order="12" place="12" resultid="42221" />
                    <RANKING order="13" place="12" resultid="43470" />
                    <RANKING order="14" place="14" resultid="43388" />
                    <RANKING order="15" place="15" resultid="42091" />
                    <RANKING order="16" place="16" resultid="42670" />
                    <RANKING order="17" place="17" resultid="43004" />
                    <RANKING order="18" place="18" resultid="42491" />
                    <RANKING order="19" place="19" resultid="42799" />
                    <RANKING order="20" place="20" resultid="42435" />
                    <RANKING order="21" place="21" resultid="42486" />
                    <RANKING order="22" place="22" resultid="43177" />
                    <RANKING order="23" place="23" resultid="42816" />
                    <RANKING order="24" place="24" resultid="43676" />
                    <RANKING order="25" place="25" resultid="43655" />
                    <RANKING order="26" place="26" resultid="41636" />
                    <RANKING order="27" place="27" resultid="43921" />
                    <RANKING order="28" place="28" resultid="41879" />
                    <RANKING order="29" place="29" resultid="43367" />
                    <RANKING order="30" place="30" resultid="43814" />
                    <RANKING order="31" place="31" resultid="43606" />
                    <RANKING order="32" place="32" resultid="42377" />
                    <RANKING order="33" place="33" resultid="42729" />
                    <RANKING order="34" place="34" resultid="43701" />
                    <RANKING order="35" place="35" resultid="43260" />
                    <RANKING order="36" place="36" resultid="42472" />
                    <RANKING order="37" place="37" resultid="42481" />
                    <RANKING order="38" place="38" resultid="42687" />
                    <RANKING order="39" place="39" resultid="43797" />
                    <RANKING order="40" place="40" resultid="42965" />
                    <RANKING order="41" place="41" resultid="43787" />
                    <RANKING order="42" place="42" resultid="43890" />
                    <RANKING order="43" place="43" resultid="44010" />
                    <RANKING order="44" place="44" resultid="41720" />
                    <RANKING order="45" place="45" resultid="41840" />
                    <RANKING order="46" place="46" resultid="41688" />
                    <RANKING order="47" place="47" resultid="43517" />
                    <RANKING order="48" place="48" resultid="42869" />
                    <RANKING order="49" place="49" resultid="42215" />
                    <RANKING order="50" place="50" resultid="42249" />
                    <RANKING order="51" place="51" resultid="44022" />
                    <RANKING order="52" place="52" resultid="43706" />
                    <RANKING order="53" place="53" resultid="42118" />
                    <RANKING order="54" place="54" resultid="42056" />
                    <RANKING order="55" place="55" resultid="43380" />
                    <RANKING order="56" place="56" resultid="42958" />
                    <RANKING order="57" place="57" resultid="43927" />
                    <RANKING order="58" place="58" resultid="43006" />
                    <RANKING order="59" place="59" resultid="41953" />
                    <RANKING order="60" place="60" resultid="43992" />
                    <RANKING order="61" place="61" resultid="43286" />
                    <RANKING order="62" place="62" resultid="43553" />
                    <RANKING order="63" place="63" resultid="43165" />
                    <RANKING order="64" place="64" resultid="43688" />
                    <RANKING order="65" place="65" resultid="42723" />
                    <RANKING order="66" place="66" resultid="43982" />
                    <RANKING order="67" place="67" resultid="41649" />
                    <RANKING order="68" place="68" resultid="43060" />
                    <RANKING order="69" place="69" resultid="41682" />
                    <RANKING order="70" place="70" resultid="42831" />
                    <RANKING order="71" place="71" resultid="44026" />
                    <RANKING order="72" place="72" resultid="43593" />
                    <RANKING order="73" place="73" resultid="43734" />
                    <RANKING order="74" place="74" resultid="43035" />
                    <RANKING order="75" place="75" resultid="43913" />
                    <RANKING order="76" place="76" resultid="43671" />
                    <RANKING order="77" place="77" resultid="43725" />
                    <RANKING order="78" place="78" resultid="42367" />
                    <RANKING order="79" place="79" resultid="42148" />
                    <RANKING order="80" place="80" resultid="41753" />
                    <RANKING order="81" place="81" resultid="42805" />
                    <RANKING order="82" place="82" resultid="44005" />
                    <RANKING order="83" place="83" resultid="41766" />
                    <RANKING order="84" place="84" resultid="43716" />
                    <RANKING order="85" place="85" resultid="41862" />
                    <RANKING order="86" place="86" resultid="42681" />
                    <RANKING order="87" place="87" resultid="43621" />
                    <RANKING order="88" place="88" resultid="42041" />
                    <RANKING order="89" place="89" resultid="43395" />
                    <RANKING order="90" place="90" resultid="43731" />
                    <RANKING order="91" place="91" resultid="41656" />
                    <RANKING order="92" place="92" resultid="43073" />
                    <RANKING order="93" place="93" resultid="42753" />
                    <RANKING order="94" place="94" resultid="43023" />
                    <RANKING order="95" place="95" resultid="42672" />
                    <RANKING order="96" place="96" resultid="41805" />
                    <RANKING order="97" place="97" resultid="43160" />
                    <RANKING order="98" place="98" resultid="41874" />
                    <RANKING order="99" place="99" resultid="43361" />
                    <RANKING order="100" place="100" resultid="43497" />
                    <RANKING order="101" place="101" resultid="42130" />
                    <RANKING order="102" place="102" resultid="43155" />
                    <RANKING order="103" place="103" resultid="43584" />
                    <RANKING order="104" place="104" resultid="43544" />
                    <RANKING order="105" place="105" resultid="41680" />
                    <RANKING order="106" place="106" resultid="42404" />
                    <RANKING order="107" place="-1" resultid="41925" />
                    <RANKING order="108" place="-1" resultid="43567" />
                    <RANKING order="109" place="-1" resultid="41532" />
                    <RANKING order="110" place="-1" resultid="41714" />
                    <RANKING order="111" place="-1" resultid="41729" />
                    <RANKING order="112" place="-1" resultid="41826" />
                    <RANKING order="113" place="-1" resultid="42026" />
                    <RANKING order="114" place="-1" resultid="42336" />
                    <RANKING order="115" place="-1" resultid="42343" />
                    <RANKING order="116" place="-1" resultid="42348" />
                    <RANKING order="117" place="-1" resultid="42425" />
                    <RANKING order="118" place="-1" resultid="42497" />
                    <RANKING order="119" place="-1" resultid="42792" />
                    <RANKING order="120" place="-1" resultid="43002" />
                    <RANKING order="121" place="-1" resultid="43146" />
                    <RANKING order="122" place="-1" resultid="43171" />
                    <RANKING order="123" place="-1" resultid="43270" />
                    <RANKING order="124" place="-1" resultid="43383" />
                    <RANKING order="125" place="-1" resultid="43511" />
                    <RANKING order="126" place="-1" resultid="43629" />
                    <RANKING order="127" place="-1" resultid="43856" />
                    <RANKING order="128" place="-1" resultid="43862" />
                    <RANKING order="129" place="-1" resultid="43999" />
                    <RANKING order="130" place="-1" resultid="41521" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45032" daytime="15:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45033" daytime="15:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="45034" daytime="15:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="45035" daytime="15:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="45036" daytime="15:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="45037" daytime="15:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="45038" daytime="15:45" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="45039" daytime="15:45" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="45040" daytime="15:45" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="45041" daytime="15:50" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="45042" daytime="15:50" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="45043" daytime="15:50" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="45044" daytime="15:55" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="45045" daytime="15:55" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="45046" daytime="16:00" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="45047" daytime="16:00" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="45048" daytime="16:00" number="17" order="17" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2430" daytime="16:05" gender="F" number="30" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45479" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42334" />
                    <RANKING order="2" place="2" resultid="42186" />
                    <RANKING order="3" place="3" resultid="43669" />
                    <RANKING order="4" place="4" resultid="42786" />
                    <RANKING order="5" place="5" resultid="42997" />
                    <RANKING order="6" place="6" resultid="42456" />
                    <RANKING order="7" place="7" resultid="42740" />
                    <RANKING order="8" place="8" resultid="43623" />
                    <RANKING order="9" place="9" resultid="42359" />
                    <RANKING order="10" place="10" resultid="42353" />
                    <RANKING order="11" place="11" resultid="42346" />
                    <RANKING order="12" place="12" resultid="42160" />
                    <RANKING order="13" place="13" resultid="43010" />
                    <RANKING order="14" place="-1" resultid="42503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45480" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42203" />
                    <RANKING order="2" place="2" resultid="43971" />
                    <RANKING order="3" place="3" resultid="43776" />
                    <RANKING order="4" place="4" resultid="43639" />
                    <RANKING order="5" place="5" resultid="42080" />
                    <RANKING order="6" place="6" resultid="43635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45481" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43415" />
                    <RANKING order="2" place="2" resultid="43781" />
                    <RANKING order="3" place="3" resultid="42239" />
                    <RANKING order="4" place="-1" resultid="42446" />
                    <RANKING order="5" place="-1" resultid="41526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45482" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42734" />
                    <RANKING order="2" place="2" resultid="42163" />
                    <RANKING order="3" place="3" resultid="43274" />
                    <RANKING order="4" place="4" resultid="42510" />
                    <RANKING order="5" place="5" resultid="42853" />
                    <RANKING order="6" place="6" resultid="41550" />
                    <RANKING order="7" place="7" resultid="42727" />
                    <RANKING order="8" place="8" resultid="41624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45483" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42085" />
                    <RANKING order="2" place="2" resultid="42124" />
                    <RANKING order="3" place="3" resultid="43873" />
                    <RANKING order="4" place="4" resultid="41973" />
                    <RANKING order="5" place="5" resultid="41947" />
                    <RANKING order="6" place="6" resultid="42717" />
                    <RANKING order="7" place="7" resultid="41817" />
                    <RANKING order="8" place="-1" resultid="41942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45484" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43304" />
                    <RANKING order="2" place="2" resultid="43682" />
                    <RANKING order="3" place="3" resultid="43754" />
                    <RANKING order="4" place="4" resultid="42244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45485" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42142" />
                    <RANKING order="2" place="2" resultid="42074" />
                    <RANKING order="3" place="3" resultid="43439" />
                    <RANKING order="4" place="4" resultid="41855" />
                    <RANKING order="5" place="5" resultid="43977" />
                    <RANKING order="6" place="6" resultid="43749" />
                    <RANKING order="7" place="7" resultid="43759" />
                    <RANKING order="8" place="8" resultid="43940" />
                    <RANKING order="9" place="9" resultid="42693" />
                    <RANKING order="10" place="10" resultid="41759" />
                    <RANKING order="11" place="11" resultid="43481" />
                    <RANKING order="12" place="12" resultid="42826" />
                    <RANKING order="13" place="13" resultid="43652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45486" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41917" />
                    <RANKING order="2" place="2" resultid="41890" />
                    <RANKING order="3" place="3" resultid="43645" />
                    <RANKING order="4" place="4" resultid="43141" />
                    <RANKING order="5" place="-1" resultid="43573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45487" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41884" />
                    <RANKING order="2" place="-1" resultid="43538" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45488" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41822" />
                    <RANKING order="2" place="2" resultid="43229" />
                    <RANKING order="3" place="-1" resultid="41708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45489" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45490" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45491" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45492" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45493" agemax="-1" agemin="-1" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42334" />
                    <RANKING order="2" place="2" resultid="42186" />
                    <RANKING order="3" place="3" resultid="43669" />
                    <RANKING order="4" place="4" resultid="42786" />
                    <RANKING order="5" place="5" resultid="42997" />
                    <RANKING order="6" place="6" resultid="43415" />
                    <RANKING order="7" place="7" resultid="42456" />
                    <RANKING order="8" place="8" resultid="42085" />
                    <RANKING order="9" place="9" resultid="42740" />
                    <RANKING order="10" place="10" resultid="43623" />
                    <RANKING order="11" place="11" resultid="42359" />
                    <RANKING order="12" place="12" resultid="42124" />
                    <RANKING order="13" place="13" resultid="42203" />
                    <RANKING order="14" place="14" resultid="43971" />
                    <RANKING order="15" place="15" resultid="43776" />
                    <RANKING order="16" place="16" resultid="42353" />
                    <RANKING order="17" place="17" resultid="43639" />
                    <RANKING order="18" place="18" resultid="43304" />
                    <RANKING order="19" place="19" resultid="42346" />
                    <RANKING order="20" place="20" resultid="42142" />
                    <RANKING order="21" place="21" resultid="42734" />
                    <RANKING order="22" place="22" resultid="43873" />
                    <RANKING order="23" place="23" resultid="41973" />
                    <RANKING order="24" place="24" resultid="42080" />
                    <RANKING order="25" place="25" resultid="42160" />
                    <RANKING order="26" place="25" resultid="43781" />
                    <RANKING order="27" place="27" resultid="42074" />
                    <RANKING order="28" place="28" resultid="43010" />
                    <RANKING order="29" place="29" resultid="42163" />
                    <RANKING order="30" place="30" resultid="43274" />
                    <RANKING order="31" place="31" resultid="41917" />
                    <RANKING order="32" place="32" resultid="43635" />
                    <RANKING order="33" place="33" resultid="43439" />
                    <RANKING order="34" place="34" resultid="42510" />
                    <RANKING order="35" place="35" resultid="41855" />
                    <RANKING order="36" place="36" resultid="42853" />
                    <RANKING order="37" place="37" resultid="43977" />
                    <RANKING order="38" place="38" resultid="41550" />
                    <RANKING order="39" place="39" resultid="41947" />
                    <RANKING order="40" place="40" resultid="43682" />
                    <RANKING order="41" place="41" resultid="43749" />
                    <RANKING order="42" place="42" resultid="42717" />
                    <RANKING order="43" place="43" resultid="42239" />
                    <RANKING order="44" place="44" resultid="43754" />
                    <RANKING order="45" place="45" resultid="42727" />
                    <RANKING order="46" place="46" resultid="43759" />
                    <RANKING order="47" place="47" resultid="43940" />
                    <RANKING order="48" place="48" resultid="42693" />
                    <RANKING order="49" place="49" resultid="42244" />
                    <RANKING order="50" place="50" resultid="41759" />
                    <RANKING order="51" place="51" resultid="41884" />
                    <RANKING order="52" place="52" resultid="41624" />
                    <RANKING order="53" place="53" resultid="41890" />
                    <RANKING order="54" place="54" resultid="43481" />
                    <RANKING order="55" place="55" resultid="42826" />
                    <RANKING order="56" place="56" resultid="43652" />
                    <RANKING order="57" place="57" resultid="43645" />
                    <RANKING order="58" place="58" resultid="41817" />
                    <RANKING order="59" place="59" resultid="43141" />
                    <RANKING order="60" place="60" resultid="41822" />
                    <RANKING order="61" place="61" resultid="43229" />
                    <RANKING order="62" place="-1" resultid="41708" />
                    <RANKING order="63" place="-1" resultid="42446" />
                    <RANKING order="64" place="-1" resultid="43538" />
                    <RANKING order="65" place="-1" resultid="43573" />
                    <RANKING order="66" place="-1" resultid="41526" />
                    <RANKING order="67" place="-1" resultid="41942" />
                    <RANKING order="68" place="-1" resultid="42503" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45065" daytime="16:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45066" daytime="16:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="45067" daytime="16:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="45068" daytime="16:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="45069" daytime="16:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="45070" daytime="16:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="45071" daytime="16:15" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="45072" daytime="16:20" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="45073" daytime="16:20" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2248" daytime="16:20" gender="M" number="31" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45299" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43087" />
                    <RANKING order="2" place="2" resultid="43607" />
                    <RANKING order="3" place="3" resultid="43342" />
                    <RANKING order="4" place="-1" resultid="43603" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45300" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43633" />
                    <RANKING order="2" place="2" resultid="42020" />
                    <RANKING order="3" place="-1" resultid="42014" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45301" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43824" />
                    <RANKING order="2" place="2" resultid="43949" />
                    <RANKING order="3" place="3" resultid="42051" />
                    <RANKING order="4" place="4" resultid="42008" />
                    <RANKING order="5" place="5" resultid="43092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45302" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42991" />
                    <RANKING order="2" place="2" resultid="41912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45303" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="41969" />
                    <RANKING order="2" place="2" resultid="41811" />
                    <RANKING order="3" place="3" resultid="41741" />
                    <RANKING order="4" place="4" resultid="42097" />
                    <RANKING order="5" place="5" resultid="43915" />
                    <RANKING order="6" place="6" resultid="43726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45304" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43318" />
                    <RANKING order="2" place="2" resultid="42478" />
                    <RANKING order="3" place="3" resultid="43261" />
                    <RANKING order="4" place="4" resultid="42183" />
                    <RANKING order="5" place="5" resultid="43841" />
                    <RANKING order="6" place="-1" resultid="42113" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45305" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43348" />
                    <RANKING order="2" place="2" resultid="42003" />
                    <RANKING order="3" place="3" resultid="41674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45306" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42976" />
                    <RANKING order="2" place="2" resultid="43523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45307" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45308" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="42747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45309" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45310" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45311" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45312" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45313" agemax="94" agemin="25" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43824" />
                    <RANKING order="2" place="2" resultid="43949" />
                    <RANKING order="3" place="3" resultid="42051" />
                    <RANKING order="4" place="4" resultid="42991" />
                    <RANKING order="5" place="5" resultid="42976" />
                    <RANKING order="6" place="6" resultid="43087" />
                    <RANKING order="7" place="7" resultid="42008" />
                    <RANKING order="8" place="8" resultid="43318" />
                    <RANKING order="9" place="9" resultid="41912" />
                    <RANKING order="10" place="10" resultid="41969" />
                    <RANKING order="11" place="11" resultid="43633" />
                    <RANKING order="12" place="12" resultid="42478" />
                    <RANKING order="13" place="13" resultid="43607" />
                    <RANKING order="14" place="14" resultid="43348" />
                    <RANKING order="15" place="15" resultid="41811" />
                    <RANKING order="16" place="16" resultid="43342" />
                    <RANKING order="17" place="17" resultid="43261" />
                    <RANKING order="18" place="18" resultid="41741" />
                    <RANKING order="19" place="19" resultid="42183" />
                    <RANKING order="20" place="20" resultid="42097" />
                    <RANKING order="21" place="21" resultid="42020" />
                    <RANKING order="22" place="22" resultid="43523" />
                    <RANKING order="23" place="23" resultid="43092" />
                    <RANKING order="24" place="24" resultid="42003" />
                    <RANKING order="25" place="25" resultid="43915" />
                    <RANKING order="26" place="26" resultid="42103" />
                    <RANKING order="27" place="27" resultid="43726" />
                    <RANKING order="28" place="28" resultid="43841" />
                    <RANKING order="29" place="29" resultid="42747" />
                    <RANKING order="30" place="30" resultid="41674" />
                    <RANKING order="31" place="-1" resultid="42014" />
                    <RANKING order="32" place="-1" resultid="42113" />
                    <RANKING order="33" place="-1" resultid="43603" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45058" daytime="16:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45059" daytime="16:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="45060" daytime="16:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="45061" daytime="16:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="45062" daytime="17:00" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2400" daytime="17:05" gender="F" number="32" order="4" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="385" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="45464" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="44036" />
                    <RANKING order="2" place="2" resultid="43298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45465" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="45466" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="45467" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43067" />
                    <RANKING order="2" place="-1" resultid="43401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45468" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43280" />
                    <RANKING order="2" place="2" resultid="43243" />
                    <RANKING order="3" place="3" resultid="43255" />
                    <RANKING order="4" place="-1" resultid="43771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45469" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43223" />
                    <RANKING order="2" place="-1" resultid="42177" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45470" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="45471" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="41705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="45472" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="45473" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="45474" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="45475" agemax="84" agemin="80" />
                <AGEGROUP agegroupid="45476" agemax="89" agemin="85" />
                <AGEGROUP agegroupid="45477" agemax="94" agemin="90" />
                <AGEGROUP agegroupid="45478" agemax="-1" agemin="-1" name="Absoluto">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="43280" />
                    <RANKING order="2" place="2" resultid="43067" />
                    <RANKING order="3" place="3" resultid="43223" />
                    <RANKING order="4" place="4" resultid="44036" />
                    <RANKING order="5" place="5" resultid="43298" />
                    <RANKING order="6" place="6" resultid="43243" />
                    <RANKING order="7" place="7" resultid="43255" />
                    <RANKING order="8" place="-1" resultid="41705" />
                    <RANKING order="9" place="-1" resultid="42177" />
                    <RANKING order="10" place="-1" resultid="43401" />
                    <RANKING order="11" place="-1" resultid="43771" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="45063" daytime="17:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="45064" daytime="17:15" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="SCA" nation="POR" region="ANCNP" clubid="43011" swrid="73233" name="Sporting Clube de Aveiro" shortname="Sporting de Aveiro">
          <ATHLETES>
            <ATHLETE firstname="Hugo Alexandre" lastname="Borrego" birthdate="1972-11-22" gender="M" nation="POR" license="205001" swrid="5220481" athleteid="43030">
              <RESULTS>
                <RESULT comment="701 - Mais de uma pernada de golfinho durante a braçada submarina - SW 7.1" eventid="2188" reactiontime="+111" status="DSQ" swimtime="00:00:51.22" resultid="43031" heatid="44942" lane="3" entrytime="00:00:45.69" entrycourse="LCM" />
                <RESULT eventid="2415" points="220" reactiontime="+118" swimtime="00:01:32.43" resultid="43032" heatid="45107" lane="8" entrytime="00:01:26.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="160" swimtime="00:00:52.95" resultid="43033" heatid="45016" lane="2" entrytime="00:00:52.31" entrycourse="LCM" />
                <RESULT eventid="2445" points="170" reactiontime="+113" swimtime="00:02:04.32" resultid="43034" heatid="44992" lane="4" entrytime="00:01:54.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="349" reactiontime="+105" swimtime="00:00:35.31" resultid="43035" heatid="45039" lane="8" entrytime="00:00:33.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jorge Vieira" lastname="Ribeiro" birthdate="1964-03-13" gender="M" nation="POR" license="128894" swrid="4939020" athleteid="43055">
              <RESULTS>
                <RESULT eventid="1058" points="343" swimtime="00:13:29.73" resultid="43056" heatid="45082" lane="3" entrytime="00:13:35.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.14" />
                    <SPLIT distance="200" swimtime="00:03:18.30" />
                    <SPLIT distance="300" swimtime="00:05:01.17" />
                    <SPLIT distance="400" swimtime="00:06:43.86" />
                    <SPLIT distance="500" swimtime="00:08:26.58" />
                    <SPLIT distance="600" swimtime="00:10:09.30" />
                    <SPLIT distance="700" swimtime="00:11:51.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2537" points="351" reactiontime="+116" swimtime="00:01:36.78" resultid="43057" heatid="44886" lane="8" entrytime="00:01:40.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.78" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="604 - Durante o percurso perdeu a posição dorsal - SW 6.2" eventid="2218" reactiontime="+95" status="DSQ" swimtime="00:03:29.73" resultid="43058" heatid="44918" lane="6" entrytime="00:03:45.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.74" />
                    <SPLIT distance="100" swimtime="00:01:41.87" />
                    <SPLIT distance="150" swimtime="00:02:36.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="400" reactiontime="+85" swimtime="00:00:42.49" resultid="43059" heatid="45018" lane="2" entrytime="00:00:43.00" entrycourse="LCM" />
                <RESULT eventid="2652" points="486" reactiontime="+112" swimtime="00:00:33.83" resultid="43060" heatid="45038" lane="3" entrytime="00:00:34.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Goncalves" lastname="Santos" birthdate="1954-03-31" gender="M" nation="POR" license="133236" swrid="5083883" athleteid="43018">
              <RESULTS>
                <RESULT eventid="2682" points="237" reactiontime="+115" swimtime="00:00:49.33" resultid="43019" heatid="44893" lane="6" entrytime="00:00:52.38" entrycourse="LCM" />
                <RESULT eventid="2323" points="164" reactiontime="+116" swimtime="00:02:13.49" resultid="43020" heatid="44925" lane="3" entrytime="00:02:06.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="251" reactiontime="+110" swimtime="00:01:39.50" resultid="43021" heatid="45105" lane="8" entrytime="00:01:38.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" points="145" reactiontime="+112" swimtime="00:05:22.33" resultid="43022" heatid="45028" lane="6" entrytime="00:05:15.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.68" />
                    <SPLIT distance="100" swimtime="00:02:33.17" />
                    <SPLIT distance="150" swimtime="00:04:05.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="315" reactiontime="+107" swimtime="00:00:41.67" resultid="43023" heatid="45035" lane="2" entrytime="00:00:40.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Maria" lastname="Martins" birthdate="1979-10-26" gender="F" nation="POR" license="123246" swrid="4756632" athleteid="43042">
              <RESULTS>
                <RESULT eventid="1060" points="222" swimtime="00:16:09.74" resultid="43043" heatid="45076" lane="8" entrytime="00:15:53.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:57.12" />
                    <SPLIT distance="200" swimtime="00:04:01.70" />
                    <SPLIT distance="300" swimtime="00:06:05.04" />
                    <SPLIT distance="400" swimtime="00:08:08.55" />
                    <SPLIT distance="500" swimtime="00:10:11.41" />
                    <SPLIT distance="600" swimtime="00:12:14.06" />
                    <SPLIT distance="700" swimtime="00:14:15.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2173" points="325" swimtime="00:04:07.00" resultid="43044" heatid="45088" lane="8" entrytime="00:04:07.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.25" />
                    <SPLIT distance="100" swimtime="00:02:00.36" />
                    <SPLIT distance="150" swimtime="00:03:04.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2203" points="201" reactiontime="+106" swimtime="00:01:59.58" resultid="43045" heatid="44881" lane="7" entrytime="00:01:56.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2308" points="213" reactiontime="+118" swimtime="00:04:17.81" resultid="43046" heatid="44914" lane="1" entrytime="00:04:04.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.19" />
                    <SPLIT distance="100" swimtime="00:02:11.40" />
                    <SPLIT distance="150" swimtime="00:03:17.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="253" reactiontime="+106" swimtime="00:03:59.32" resultid="43047" heatid="44971" lane="5" entrytime="00:04:07.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.63" />
                    <SPLIT distance="100" swimtime="00:02:06.32" />
                    <SPLIT distance="150" swimtime="00:03:08.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eliana Marta" lastname="Castro" birthdate="1970-12-02" gender="F" nation="POR" license="214221" athleteid="43053">
              <RESULTS>
                <RESULT eventid="2308" points="196" reactiontime="+183" swimtime="00:04:42.39" resultid="43054" heatid="44913" lane="2" entrytime="00:04:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.39" />
                    <SPLIT distance="100" swimtime="00:02:18.93" />
                    <SPLIT distance="150" swimtime="00:03:33.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Alexandre" lastname="Raposo" birthdate="1955-06-18" gender="M" nation="POR" license="131484" swrid="5027372" athleteid="43024">
              <RESULTS>
                <RESULT eventid="2537" points="204" reactiontime="+75" swimtime="00:02:05.34" resultid="43025" heatid="44885" lane="7" entrytime="00:01:58.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="210" reactiontime="+82" swimtime="00:04:30.43" resultid="43026" heatid="44916" lane="4" entrytime="00:04:36.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.14" />
                    <SPLIT distance="100" swimtime="00:02:13.70" />
                    <SPLIT distance="150" swimtime="00:03:22.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="247" reactiontime="+100" swimtime="00:01:40.05" resultid="43027" heatid="45104" lane="4" entrytime="00:01:41.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="275" reactiontime="+99" swimtime="00:08:03.23" resultid="43028" heatid="45125" lane="1" entrytime="00:08:13.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.63" />
                    <SPLIT distance="100" swimtime="00:01:55.29" />
                    <SPLIT distance="150" swimtime="00:02:57.80" />
                    <SPLIT distance="200" swimtime="00:04:01.33" />
                    <SPLIT distance="250" swimtime="00:05:03.37" />
                    <SPLIT distance="300" swimtime="00:06:05.18" />
                    <SPLIT distance="350" swimtime="00:07:05.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="205" reactiontime="+87" swimtime="00:00:56.75" resultid="43029" heatid="45016" lane="7" entrytime="00:00:52.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Claudia Baptista" lastname="Domingues" birthdate="1977-05-04" gender="F" nation="POR" license="203924" swrid="4003289" athleteid="43036">
              <RESULTS>
                <RESULT eventid="2338" points="553" reactiontime="+86" swimtime="00:00:35.74" resultid="43037" heatid="44892" lane="1" entrytime="00:00:35.66" entrycourse="LCM" />
                <RESULT eventid="2278" points="403" reactiontime="+97" swimtime="00:02:58.15" resultid="43038" heatid="44904" lane="5" entrytime="00:02:51.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                    <SPLIT distance="100" swimtime="00:01:23.41" />
                    <SPLIT distance="150" swimtime="00:02:11.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="509" reactiontime="+88" swimtime="00:01:15.50" resultid="43039" heatid="44956" lane="6" entrytime="00:01:14.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="478" reactiontime="+96" swimtime="00:03:13.65" resultid="43040" heatid="44972" lane="5" entrytime="00:03:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:01:28.36" />
                    <SPLIT distance="150" swimtime="00:02:27.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="453" reactiontime="+112" swimtime="00:00:41.21" resultid="43041" heatid="45026" lane="8" entrytime="00:00:41.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel Castro" lastname="Trigo" birthdate="1965-11-25" gender="M" nation="POR" license="120704" swrid="4652887" athleteid="43012">
              <RESULTS>
                <RESULT eventid="1058" points="267" swimtime="00:14:39.99" resultid="43013" heatid="45081" lane="6" entrytime="00:14:14.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.02" />
                    <SPLIT distance="200" swimtime="00:03:33.46" />
                    <SPLIT distance="300" swimtime="00:05:27.27" />
                    <SPLIT distance="400" swimtime="00:07:20.49" />
                    <SPLIT distance="500" swimtime="00:09:13.44" />
                    <SPLIT distance="600" swimtime="00:11:04.07" />
                    <SPLIT distance="700" swimtime="00:12:54.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2622" points="340" reactiontime="+103" swimtime="00:03:54.08" resultid="43014" heatid="44875" lane="6" entrytime="00:03:41.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.85" />
                    <SPLIT distance="100" swimtime="00:01:55.42" />
                    <SPLIT distance="150" swimtime="00:02:55.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="218" reactiontime="+88" swimtime="00:04:10.61" resultid="43015" heatid="44918" lane="1" entrytime="00:03:50.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.25" />
                    <SPLIT distance="100" swimtime="00:02:05.58" />
                    <SPLIT distance="150" swimtime="00:03:09.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="304" reactiontime="+101" swimtime="00:00:46.14" resultid="43016" heatid="44943" lane="8" entrytime="00:00:45.08" entrycourse="LCM" />
                <RESULT eventid="2385" points="240" reactiontime="+119" swimtime="00:04:06.38" resultid="43017" heatid="44976" lane="3" entrytime="00:03:43.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.47" />
                    <SPLIT distance="100" swimtime="00:02:01.05" />
                    <SPLIT distance="150" swimtime="00:03:12.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Celso Abreu" lastname="Fernandes" birthdate="1967-11-06" gender="M" nation="POR" license="213521" swrid="5450760" athleteid="43048">
              <RESULTS>
                <RESULT eventid="2537" points="146" reactiontime="+131" swimtime="00:02:05.06" resultid="43049" heatid="44884" lane="5" entrytime="00:02:10.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="221" reactiontime="+117" swimtime="00:03:30.27" resultid="43050" heatid="45091" lane="5" entrytime="00:03:20.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.38" />
                    <SPLIT distance="100" swimtime="00:01:41.08" />
                    <SPLIT distance="150" swimtime="00:02:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="151" reactiontime="+109" swimtime="00:00:58.36" resultid="43051" heatid="44938" lane="5" entrytime="00:01:01.16" entrycourse="LCM" />
                <RESULT eventid="2445" points="199" reactiontime="+121" swimtime="00:02:04.06" resultid="43052" heatid="44991" lane="3" entrytime="00:02:09.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CCLAMAS" nation="POR" region="ANNP" clubid="42354" swrid="68108" name="Clube Colegio de Lamas" shortname="Colegio SMLamas">
          <ATHLETES>
            <ATHLETE firstname="Diana Maria" lastname="Espinheira" birthdate="1992-02-11" gender="F" nation="POR" license="103996" swrid="4123303" athleteid="42360">
              <RESULTS>
                <RESULT eventid="2607" points="403" reactiontime="+89" swimtime="00:00:44.20" resultid="42361" heatid="45102" lane="1" entrytime="00:00:44.13" entrycourse="LCM" />
                <RESULT eventid="2460" points="402" reactiontime="+90" swimtime="00:01:38.00" resultid="42362" heatid="45122" lane="6" entrytime="00:01:38.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alberto Nuno" lastname="Espinheiro" birthdate="1962-08-11" gender="M" nation="POR" license="106811" swrid="4372683" athleteid="42363">
              <RESULTS>
                <RESULT eventid="2188" points="346" reactiontime="+88" swimtime="00:00:44.21" resultid="42364" heatid="44944" lane="4" entrytime="00:00:43.24" entrycourse="LCM" />
                <RESULT eventid="2415" points="332" reactiontime="+92" swimtime="00:01:26.77" resultid="42365" heatid="45106" lane="1" entrytime="00:01:28.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="360" reactiontime="+86" swimtime="00:01:42.07" resultid="42366" heatid="44995" lane="6" entrytime="00:01:37.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="399" reactiontime="+86" swimtime="00:00:36.14" resultid="42367" heatid="45036" lane="8" entrytime="00:00:38.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Lucia" lastname="Castro" birthdate="1992-12-18" gender="F" nation="POR" license="102795" swrid="4123671" athleteid="42355">
              <RESULTS>
                <RESULT eventid="2173" points="563" swimtime="00:03:08.68" resultid="42356" heatid="45089" lane="3" entrytime="00:03:11.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="100" swimtime="00:01:30.93" />
                    <SPLIT distance="150" swimtime="00:02:19.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="632" reactiontime="+86" swimtime="00:00:38.04" resultid="42357" heatid="45103" lane="6" entrytime="00:00:37.98" entrycourse="LCM" />
                <RESULT eventid="2460" points="637" reactiontime="+82" swimtime="00:01:24.10" resultid="42358" heatid="45123" lane="6" entrytime="00:01:28.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="582" reactiontime="+82" swimtime="00:00:31.26" resultid="42359" heatid="45073" lane="1" entrytime="00:00:30.36" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur Sousa" lastname="Ferreira" birthdate="1993-02-21" gender="M" nation="POR" license="108511" swrid="4345551" athleteid="42368">
              <RESULTS>
                <RESULT eventid="2507" points="540" reactiontime="+76" swimtime="00:02:21.38" resultid="42369" heatid="45095" lane="3" entrytime="00:02:19.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:07.60" />
                    <SPLIT distance="150" swimtime="00:01:43.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="589" reactiontime="+81" swimtime="00:01:01.68" resultid="42370" heatid="45115" lane="8" entrytime="00:01:00.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="553" reactiontime="+92" swimtime="00:05:05.62" resultid="42371" heatid="45131" lane="1" entrytime="00:05:07.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:09.31" />
                    <SPLIT distance="150" swimtime="00:01:47.49" />
                    <SPLIT distance="200" swimtime="00:02:26.64" />
                    <SPLIT distance="250" swimtime="00:03:06.26" />
                    <SPLIT distance="300" swimtime="00:03:46.23" />
                    <SPLIT distance="350" swimtime="00:04:25.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="595" reactiontime="+75" swimtime="00:00:27.52" resultid="42372" heatid="45046" lane="2" entrytime="00:00:27.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme Araujo" lastname="Soares" birthdate="1993-11-02" gender="M" nation="POR" license="111295" swrid="4397502" athleteid="42373">
              <RESULTS>
                <RESULT eventid="2682" points="561" reactiontime="+73" swimtime="00:00:30.38" resultid="42374" heatid="44900" lane="1" entrytime="00:00:29.70" entrycourse="LCM" />
                <RESULT eventid="2323" points="574" reactiontime="+66" swimtime="00:01:08.40" resultid="42375" heatid="44928" lane="6" entrytime="00:01:10.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="450" reactiontime="+75" swimtime="00:00:34.94" resultid="42376" heatid="45020" lane="8" entrytime="00:00:35.61" entrycourse="SCM" />
                <RESULT eventid="2652" points="514" reactiontime="+65" swimtime="00:00:28.90" resultid="42377" heatid="45044" lane="3" entrytime="00:00:28.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CCDSERTA" nation="POR" region="ANIC" clubid="41538" swrid="85400" name="CCD Pess. Camara Munic. da Serta" shortname="CCDSerta">
          <ATHLETES>
            <ATHLETE firstname="Ingrid Bernadette" lastname="Thuillier" birthdate="1981-05-21" gender="F" nation="FRA" license="212625" swrid="5429047" athleteid="41545">
              <RESULTS>
                <RESULT eventid="2278" points="266" reactiontime="+109" swimtime="00:03:24.56" resultid="41546" heatid="44903" lane="2" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.88" />
                    <SPLIT distance="100" swimtime="00:01:40.45" />
                    <SPLIT distance="150" swimtime="00:02:35.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="437" reactiontime="+100" swimtime="00:00:46.05" resultid="41547" heatid="45099" lane="7" entrytime="00:00:52.51" entrycourse="SCM" />
                <RESULT eventid="2637" points="290" reactiontime="+88" swimtime="00:01:31.10" resultid="41548" heatid="44954" lane="6" entrytime="00:01:31.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="316" reactiontime="+82" swimtime="00:01:52.66" resultid="41549" heatid="45120" lane="6" entrytime="00:01:51.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="352" reactiontime="+86" swimtime="00:00:38.87" resultid="41550" heatid="45067" lane="3" entrytime="00:00:45.10" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laurelin Lucinda" lastname="Molen" birthdate="1987-12-22" gender="F" nation="NED" license="210456" swrid="5361375" athleteid="41539">
              <RESULTS>
                <RESULT eventid="1060" points="330" swimtime="00:13:36.86" resultid="41540" heatid="45077" lane="5" entrytime="00:13:20.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.61" />
                    <SPLIT distance="200" swimtime="00:03:16.46" />
                    <SPLIT distance="300" swimtime="00:05:00.94" />
                    <SPLIT distance="400" swimtime="00:06:45.37" />
                    <SPLIT distance="500" swimtime="00:08:30.20" />
                    <SPLIT distance="600" swimtime="00:10:14.47" />
                    <SPLIT distance="700" swimtime="00:11:56.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2173" points="400" swimtime="00:03:36.15" resultid="41541" heatid="45089" lane="2" entrytime="00:03:30.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.98" />
                    <SPLIT distance="100" swimtime="00:01:43.53" />
                    <SPLIT distance="150" swimtime="00:02:40.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2278" points="285" reactiontime="+91" swimtime="00:03:13.65" resultid="41542" heatid="44904" lane="1" entrytime="00:03:07.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.56" />
                    <SPLIT distance="100" swimtime="00:01:30.70" />
                    <SPLIT distance="150" swimtime="00:02:22.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="337" reactiontime="+90" swimtime="00:06:32.84" resultid="41543" heatid="45012" lane="6" entrytime="00:06:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                    <SPLIT distance="100" swimtime="00:01:30.30" />
                    <SPLIT distance="150" swimtime="00:02:19.45" />
                    <SPLIT distance="200" swimtime="00:03:10.09" />
                    <SPLIT distance="250" swimtime="00:04:00.91" />
                    <SPLIT distance="300" swimtime="00:04:51.72" />
                    <SPLIT distance="350" swimtime="00:05:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="364" reactiontime="+96" swimtime="00:01:40.76" resultid="41544" heatid="45122" lane="3" entrytime="00:01:37.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ANE" nation="POR" region="ANL" clubid="41527" swrid="73259" name="CCD Associacao de Nadadores dos Estoris" shortname="Nadadores dos Estoris">
          <ATHLETES>
            <ATHLETE firstname="Ruben Tiago" lastname="Perdigoto" birthdate="1989-10-04" gender="M" nation="POR" license="205088" swrid="5231594" athleteid="41528">
              <RESULTS>
                <RESULT eventid="2682" status="DNS" swimtime="00:00:00.00" resultid="41529" heatid="44899" lane="4" entrytime="00:00:29.90" />
                <RESULT eventid="2323" status="DNS" swimtime="00:00:00.00" resultid="41530" heatid="44929" lane="8" entrytime="00:01:09.00" />
                <RESULT eventid="2415" status="DNS" swimtime="00:00:00.00" resultid="41531" heatid="45115" lane="2" entrytime="00:01:00.00" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="41532" heatid="45047" lane="6" entrytime="00:00:26.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ralf Pinto" lastname="Soares" birthdate="1964-08-02" gender="M" nation="POR" license="26786" swrid="4575903" athleteid="41533">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="41534" heatid="45082" lane="7" entrytime="00:13:45.00" />
                <RESULT eventid="2622" status="DNS" swimtime="00:00:00.00" resultid="41535" heatid="44877" lane="2" entrytime="00:03:19.50" />
                <RESULT eventid="2507" status="DNS" swimtime="00:00:00.00" resultid="41536" heatid="45093" lane="3" entrytime="00:02:45.00" />
                <RESULT eventid="2385" status="DNS" swimtime="00:00:00.00" resultid="41537" heatid="44978" lane="6" entrytime="00:03:10.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GCST" nation="POR" region="ANNP" clubid="42870" swrid="68074" name="Ginasio Clube de Santo Tirso" shortname="Ginasio Santo Tirso">
          <ATHLETES>
            <ATHLETE firstname="Delfina Maria" lastname="Martins" birthdate="1966-11-22" gender="F" nation="POR" license="117387" swrid="4496950" athleteid="43648">
              <RESULTS>
                <RESULT eventid="1060" points="163" swimtime="00:18:25.85" resultid="43649" heatid="45075" lane="2" entrytime="00:17:18.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:10.33" />
                    <SPLIT distance="200" swimtime="00:04:27.84" />
                    <SPLIT distance="300" swimtime="00:06:47.18" />
                    <SPLIT distance="400" swimtime="00:09:07.01" />
                    <SPLIT distance="500" swimtime="00:11:26.58" />
                    <SPLIT distance="600" swimtime="00:13:46.42" />
                    <SPLIT distance="700" swimtime="00:16:07.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2278" points="152" reactiontime="+131" swimtime="00:04:21.44" resultid="43650" heatid="44902" lane="2" entrytime="00:04:10.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.53" />
                    <SPLIT distance="100" swimtime="00:02:07.04" />
                    <SPLIT distance="150" swimtime="00:03:14.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="144" reactiontime="+131" swimtime="00:02:01.43" resultid="43651" heatid="44952" lane="6" entrytime="00:01:58.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="161" reactiontime="+131" swimtime="00:00:54.36" resultid="43652" heatid="45066" lane="5" entrytime="00:00:52.51" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariana Dias" lastname="Almeida" birthdate="1993-09-12" gender="F" nation="POR" license="22405" swrid="4074209" athleteid="43622">
              <RESULTS>
                <RESULT eventid="2430" points="588" reactiontime="+76" swimtime="00:00:31.14" resultid="43623" heatid="45073" lane="2" entrytime="00:00:30.06" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Eduardo" lastname="Afonso" birthdate="1965-11-07" gender="M" nation="POR" license="207922" swrid="5032171" athleteid="43618">
              <RESULTS>
                <RESULT comment="815 - Na chegada tocou com uma mão - SW 8.4" eventid="2682" reactiontime="+85" status="DSQ" swimtime="00:00:45.13" resultid="43619" heatid="44894" lane="1" entrytime="00:00:46.20" entrycourse="SCM" />
                <RESULT eventid="2188" points="361" reactiontime="+84" swimtime="00:00:43.60" resultid="43620" heatid="44945" lane="1" entrytime="00:00:43.18" entrycourse="SCM" />
                <RESULT eventid="2652" points="323" reactiontime="+80" swimtime="00:00:38.76" resultid="43621" heatid="45035" lane="7" entrytime="00:00:40.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cristiano Rocha" lastname="Ferreira" birthdate="1973-02-17" gender="M" nation="POR" license="131837" swrid="5041323" athleteid="43627">
              <RESULTS>
                <RESULT eventid="2188" status="DNS" swimtime="00:00:00.00" resultid="43628" heatid="44940" lane="5" entrytime="00:00:50.18" entrycourse="LCM" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="43629" heatid="45036" lane="2" entrytime="00:00:37.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gracinda Maria" lastname="Machado" birthdate="1961-05-01" gender="F" nation="POR" license="117386" swrid="4496949" athleteid="43642">
              <RESULTS>
                <RESULT eventid="1060" points="229" swimtime="00:19:14.88" resultid="43643" heatid="45074" lane="1" entrytime="00:20:02.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:11.40" />
                    <SPLIT distance="200" swimtime="00:04:34.27" />
                    <SPLIT distance="300" swimtime="00:06:59.90" />
                    <SPLIT distance="400" swimtime="00:09:26.53" />
                    <SPLIT distance="500" swimtime="00:11:55.17" />
                    <SPLIT distance="600" swimtime="00:14:23.61" />
                    <SPLIT distance="700" swimtime="00:16:52.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="173" reactiontime="+108" swimtime="00:02:06.07" resultid="43644" heatid="44952" lane="1" entrytime="00:02:11.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="178" reactiontime="+106" swimtime="00:00:55.34" resultid="43645" heatid="45066" lane="2" entrytime="00:00:57.99" entrycourse="SCM" />
                <RESULT eventid="2173" points="235" swimtime="00:05:17.03" resultid="43646" heatid="45086" lane="4" entrytime="00:04:57.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.99" />
                    <SPLIT distance="100" swimtime="00:02:33.99" />
                    <SPLIT distance="150" swimtime="00:03:57.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="190" reactiontime="+107" swimtime="00:02:29.11" resultid="43647" heatid="45118" lane="3" entrytime="00:02:21.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Augusto Mariano" lastname="Soares" birthdate="1972-03-05" gender="M" nation="POR" license="117424" swrid="4496951" athleteid="43656">
              <RESULTS>
                <RESULT eventid="2293" points="95" reactiontime="+69" swimtime="00:01:03.03" resultid="43657" heatid="45015" lane="6" entrytime="00:00:56.30" entrycourse="LCM" />
                <RESULT eventid="2445" points="81" swimtime="00:02:39.19" resultid="43658" heatid="44990" lane="5" entrytime="00:02:20.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:20.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Raquel" lastname="Lirio" birthdate="1990-12-10" gender="F" nation="POR" license="15206" swrid="4074207" athleteid="43640">
              <RESULTS>
                <RESULT eventid="2233" points="338" reactiontime="+98" swimtime="00:03:26.63" resultid="43641" heatid="44972" lane="4" entrytime="00:03:18.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.89" />
                    <SPLIT distance="100" swimtime="00:01:38.77" />
                    <SPLIT distance="150" swimtime="00:02:37.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rute Sofia" lastname="Teixeira" birthdate="1990-09-10" gender="F" nation="POR" license="15202" swrid="4074211" athleteid="43659">
              <RESULTS>
                <RESULT eventid="1060" points="520" swimtime="00:11:42.51" resultid="43660" heatid="45078" lane="7" entrytime="00:12:09.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.35" />
                    <SPLIT distance="200" swimtime="00:02:50.52" />
                    <SPLIT distance="300" swimtime="00:04:20.07" />
                    <SPLIT distance="400" swimtime="00:05:50.11" />
                    <SPLIT distance="500" swimtime="00:07:19.67" />
                    <SPLIT distance="600" swimtime="00:08:49.34" />
                    <SPLIT distance="700" swimtime="00:10:16.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2338" points="652" reactiontime="+85" swimtime="00:00:32.97" resultid="43661" heatid="44892" lane="2" entrytime="00:00:33.52" entrycourse="SCM" />
                <RESULT eventid="2552" points="612" reactiontime="+93" swimtime="00:01:16.01" resultid="43662" heatid="44924" lane="7" entrytime="00:01:14.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="561" reactiontime="+89" swimtime="00:05:31.71" resultid="43663" heatid="45013" lane="7" entrytime="00:05:35.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:18.09" />
                    <SPLIT distance="150" swimtime="00:02:01.04" />
                    <SPLIT distance="200" swimtime="00:02:43.95" />
                    <SPLIT distance="250" swimtime="00:03:25.79" />
                    <SPLIT distance="300" swimtime="00:04:08.27" />
                    <SPLIT distance="350" swimtime="00:04:51.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sandra Santa" lastname="Barbara" birthdate="1975-03-22" gender="F" nation="POR" license="104504" swrid="4426885" athleteid="43624">
              <RESULTS>
                <RESULT eventid="1060" points="215" swimtime="00:16:08.05" resultid="43625" heatid="45077" lane="3" entrytime="00:13:24.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.31" />
                    <SPLIT distance="200" swimtime="00:03:32.08" />
                    <SPLIT distance="300" swimtime="00:05:36.06" />
                    <SPLIT distance="400" swimtime="00:07:41.49" />
                    <SPLIT distance="500" swimtime="00:09:49.18" />
                    <SPLIT distance="600" swimtime="00:11:56.81" />
                    <SPLIT distance="700" swimtime="00:14:02.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="394" reactiontime="+86" swimtime="00:01:49.23" resultid="43626" heatid="45122" lane="2" entrytime="00:01:38.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Rosario" lastname="Figueiredo" birthdate="1989-11-02" gender="M" nation="POR" license="131311" swrid="5019410" athleteid="43630">
              <RESULTS>
                <RESULT eventid="2507" points="402" reactiontime="+80" swimtime="00:02:36.77" resultid="43631" heatid="45095" lane="2" entrytime="00:02:25.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                    <SPLIT distance="100" swimtime="00:01:12.18" />
                    <SPLIT distance="150" swimtime="00:01:54.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="434" reactiontime="+80" swimtime="00:01:07.14" resultid="43632" heatid="45112" lane="8" entrytime="00:01:06.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="335" reactiontime="+84" swimtime="00:06:34.18" resultid="43633" heatid="45060" lane="1" entrytime="00:06:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                    <SPLIT distance="100" swimtime="00:01:31.07" />
                    <SPLIT distance="150" swimtime="00:02:22.61" />
                    <SPLIT distance="200" swimtime="00:03:16.57" />
                    <SPLIT distance="250" swimtime="00:04:10.99" />
                    <SPLIT distance="300" swimtime="00:05:05.84" />
                    <SPLIT distance="350" swimtime="00:05:52.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Joao" lastname="Jose" birthdate="1990-12-17" gender="F" nation="POR" license="15208" swrid="4575034" athleteid="43636">
              <RESULTS>
                <RESULT eventid="2637" points="365" reactiontime="+91" swimtime="00:01:21.45" resultid="43637" heatid="44956" lane="4" entrytime="00:01:12.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="398" reactiontime="+82" swimtime="00:00:42.14" resultid="43638" heatid="45025" lane="4" entrytime="00:00:41.69" entrycourse="SCM" />
                <RESULT eventid="2430" points="517" reactiontime="+91" swimtime="00:00:32.96" resultid="43639" heatid="45071" lane="4" entrytime="00:00:32.39" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena Manuel" lastname="Jose" birthdate="1990-12-17" gender="F" nation="POR" license="15205" swrid="4575033" athleteid="43634">
              <RESULTS>
                <RESULT eventid="2430" points="382" reactiontime="+93" swimtime="00:00:36.46" resultid="43635" heatid="45072" lane="1" entrytime="00:00:31.99" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno Miguel" lastname="Oliveira" birthdate="1989-05-03" gender="M" nation="POR" license="207923" swrid="5065753" athleteid="43653">
              <RESULTS>
                <RESULT eventid="2415" points="439" reactiontime="+77" swimtime="00:01:06.85" resultid="43654" heatid="45111" lane="8" entrytime="00:01:09.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="546" reactiontime="+80" swimtime="00:00:28.43" resultid="43655" heatid="45042" lane="1" entrytime="00:00:30.33" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00663" nation="ESP" region="10114" clubid="41788" swrid="67670" name="C.D. Natacion Cordoba" shortname="Natacion Cordoba">
          <ATHLETES>
            <ATHLETE firstname="Marco Antonio" lastname="Castilla Gomez" birthdate="1973-06-26" gender="M" nation="ESP" swrid="4595949" athleteid="41789">
              <RESULTS>
                <RESULT eventid="2682" points="598" reactiontime="+79" swimtime="00:00:31.51" resultid="41790" heatid="44899" lane="2" entrytime="00:00:30.51" entrycourse="LCM" />
                <RESULT eventid="2323" points="565" reactiontime="+78" swimtime="00:01:13.07" resultid="41791" heatid="44929" lane="2" entrytime="00:01:07.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" points="500" reactiontime="+103" swimtime="00:02:55.47" resultid="41792" heatid="45030" lane="2" entrytime="00:02:38.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.22" />
                    <SPLIT distance="100" swimtime="00:01:24.26" />
                    <SPLIT distance="150" swimtime="00:02:12.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CDN" nation="POR" region="ANMAD" clubid="41630" swrid="65886" name="Clube Desportivo Nacional" shortname="Desportivo Nacional">
          <ATHLETES>
            <ATHLETE firstname="Duarte Nuno" lastname="Camacho" birthdate="1969-08-05" gender="M" nation="POR" license="12435" swrid="4574503" athleteid="41631">
              <RESULTS>
                <RESULT eventid="2682" points="762" reactiontime="+76" swimtime="00:00:30.25" resultid="41632" heatid="44900" lane="7" entrytime="00:00:29.50" />
                <RESULT eventid="2507" points="729" reactiontime="+76" swimtime="00:02:21.36" resultid="41633" heatid="45095" lane="4" entrytime="00:02:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                    <SPLIT distance="100" swimtime="00:01:09.07" />
                    <SPLIT distance="150" swimtime="00:01:45.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2323" points="771" reactiontime="+86" swimtime="00:01:09.45" resultid="41634" heatid="44930" lane="8" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="602" reactiontime="+77" swimtime="00:00:35.24" resultid="41635" heatid="45020" lane="6" entrytime="00:00:34.38" />
                <RESULT eventid="2652" points="689" reactiontime="+76" swimtime="00:00:28.44" resultid="41636" heatid="45046" lane="1" entrytime="00:00:27.61" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="OC" nation="POR" region="ANDL" clubid="41643" swrid="78570" name="Obidos Criativa, EEM" shortname="Obidos Criativa">
          <ATHLETES>
            <ATHLETE firstname="Daniel Rocha" lastname="Tomas" birthdate="1983-01-27" gender="M" nation="POR" license="210528" swrid="5418282" athleteid="41644">
              <RESULTS>
                <RESULT eventid="2622" points="278" reactiontime="+93" swimtime="00:03:51.74" resultid="41645" heatid="44876" lane="7" entrytime="00:03:30.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.05" />
                    <SPLIT distance="100" swimtime="00:01:47.06" />
                    <SPLIT distance="150" swimtime="00:02:50.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="245" reactiontime="+108" swimtime="00:00:40.77" resultid="41646" heatid="44895" lane="1" entrytime="00:00:40.10" entrycourse="LCM" />
                <RESULT eventid="2415" points="275" reactiontime="+100" swimtime="00:01:19.87" resultid="41647" heatid="45107" lane="3" entrytime="00:01:22.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="237" reactiontime="+104" swimtime="00:00:43.56" resultid="41648" heatid="45018" lane="8" entrytime="00:00:43.44" />
                <RESULT eventid="2652" points="341" reactiontime="+82" swimtime="00:00:33.67" resultid="41649" heatid="45039" lane="5" entrytime="00:00:33.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LPS" nation="POR" region="ANL" clubid="41997" swrid="77058" name="BJWHF Sports Club - Lisboa PoolSharks" name.en="Lisboa PoolSharks" shortname="Lisboa PoolSharks">
          <ATHLETES>
            <ATHLETE firstname="Andre Manuel" lastname="Fernandes" birthdate="1988-08-31" gender="M" nation="POR" license="208967" swrid="4800169" athleteid="42015">
              <RESULTS>
                <RESULT eventid="2622" points="310" reactiontime="+101" swimtime="00:03:31.81" resultid="42016" heatid="44876" lane="6" entrytime="00:03:28.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.58" />
                    <SPLIT distance="100" swimtime="00:01:41.39" />
                    <SPLIT distance="150" swimtime="00:02:37.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2537" points="217" reactiontime="+84" swimtime="00:01:33.98" resultid="42017" heatid="44887" lane="7" entrytime="00:01:29.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="252" reactiontime="+82" swimtime="00:03:25.69" resultid="42018" heatid="44919" lane="6" entrytime="00:03:16.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.30" />
                    <SPLIT distance="100" swimtime="00:01:38.77" />
                    <SPLIT distance="150" swimtime="00:02:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="314" reactiontime="+101" swimtime="00:03:13.58" resultid="42019" heatid="44978" lane="1" entrytime="00:03:10.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.38" />
                    <SPLIT distance="100" swimtime="00:01:33.95" />
                    <SPLIT distance="150" swimtime="00:02:26.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="264" reactiontime="+101" swimtime="00:07:06.88" resultid="42020" heatid="45059" lane="4" entrytime="00:07:19.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.70" />
                    <SPLIT distance="100" swimtime="00:01:43.07" />
                    <SPLIT distance="150" swimtime="00:02:35.54" />
                    <SPLIT distance="200" swimtime="00:03:29.61" />
                    <SPLIT distance="250" swimtime="00:04:24.96" />
                    <SPLIT distance="300" swimtime="00:05:22.94" />
                    <SPLIT distance="350" swimtime="00:06:16.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno Miguel" lastname="Silva" birthdate="1986-09-15" gender="M" nation="POR" license="210310" swrid="5345494" athleteid="42052">
              <RESULTS>
                <RESULT eventid="2622" points="429" reactiontime="+103" swimtime="00:03:20.64" resultid="42053" heatid="44878" lane="2" entrytime="00:03:13.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.90" />
                    <SPLIT distance="100" swimtime="00:01:32.39" />
                    <SPLIT distance="150" swimtime="00:02:25.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="408" reactiontime="+99" swimtime="00:00:39.36" resultid="42054" heatid="44948" lane="3" entrytime="00:00:37.68" />
                <RESULT eventid="2445" points="411" reactiontime="+83" swimtime="00:01:29.34" resultid="42055" heatid="44997" lane="4" entrytime="00:01:25.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="383" reactiontime="+78" swimtime="00:00:32.39" resultid="42056" heatid="45040" lane="7" entrytime="00:00:32.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patricia Diogenes" lastname="Pereira" birthdate="1969-11-11" gender="F" nation="POR" license="26793" swrid="4575492" athleteid="42042">
              <RESULTS>
                <RESULT eventid="1060" points="613" swimtime="00:11:36.99" resultid="42043" heatid="45078" lane="2" entrytime="00:12:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.01" />
                    <SPLIT distance="200" swimtime="00:02:50.50" />
                    <SPLIT distance="300" swimtime="00:04:18.16" />
                    <SPLIT distance="400" swimtime="00:05:45.87" />
                    <SPLIT distance="500" swimtime="00:07:14.61" />
                    <SPLIT distance="600" swimtime="00:08:43.08" />
                    <SPLIT distance="700" swimtime="00:10:10.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2173" points="613" swimtime="00:03:35.61" resultid="42044" heatid="45088" lane="5" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.24" />
                    <SPLIT distance="100" swimtime="00:01:42.58" />
                    <SPLIT distance="150" swimtime="00:02:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2308" points="598" reactiontime="+71" swimtime="00:03:14.68" resultid="42045" heatid="44914" lane="4" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.92" />
                    <SPLIT distance="100" swimtime="00:01:36.08" />
                    <SPLIT distance="150" swimtime="00:02:26.33" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rec Nac Esc F" eventid="2233" points="651" reactiontime="+77" swimtime="00:03:02.00" resultid="42046" heatid="44973" lane="1" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:25.18" />
                    <SPLIT distance="150" swimtime="00:02:21.27" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rec Nac Esc F" eventid="2492" points="652" reactiontime="+82" swimtime="00:05:32.36" resultid="42047" heatid="45013" lane="8" entrytime="00:05:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.91" />
                    <SPLIT distance="100" swimtime="00:01:16.60" />
                    <SPLIT distance="150" swimtime="00:01:58.71" />
                    <SPLIT distance="200" swimtime="00:02:40.72" />
                    <SPLIT distance="250" swimtime="00:03:23.96" />
                    <SPLIT distance="300" swimtime="00:04:06.86" />
                    <SPLIT distance="350" swimtime="00:04:50.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Miguel" lastname="Oliveira" birthdate="1983-02-26" gender="M" nation="POR" license="100486" swrid="5260317" athleteid="42032">
              <RESULTS>
                <RESULT eventid="2323" points="225" reactiontime="+111" swimtime="00:01:35.60" resultid="42033" heatid="44926" lane="5" entrytime="00:01:30.82">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="308" reactiontime="+112" swimtime="00:01:38.32" resultid="42034" heatid="44996" lane="8" entrytime="00:01:35.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="281" reactiontime="+98" swimtime="00:06:31.25" resultid="42035" heatid="45128" lane="6" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                    <SPLIT distance="100" swimtime="00:01:26.16" />
                    <SPLIT distance="150" swimtime="00:02:15.37" />
                    <SPLIT distance="200" swimtime="00:03:05.66" />
                    <SPLIT distance="250" swimtime="00:03:57.25" />
                    <SPLIT distance="300" swimtime="00:04:49.41" />
                    <SPLIT distance="350" swimtime="00:05:41.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alvaro Miguel" lastname="Cardoso" birthdate="1984-01-29" gender="M" nation="POR" license="124917" swrid="4004843" athleteid="42004">
              <RESULTS>
                <RESULT eventid="2218" points="497" reactiontime="+92" swimtime="00:02:48.13" resultid="42005" heatid="44921" lane="8" entrytime="00:02:46.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.62" />
                    <SPLIT distance="100" swimtime="00:01:20.88" />
                    <SPLIT distance="150" swimtime="00:02:04.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="517" reactiontime="+86" swimtime="00:05:19.51" resultid="42006" heatid="45130" lane="3" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:01:12.02" />
                    <SPLIT distance="150" swimtime="00:01:51.72" />
                    <SPLIT distance="200" swimtime="00:02:33.03" />
                    <SPLIT distance="250" swimtime="00:03:13.83" />
                    <SPLIT distance="300" swimtime="00:03:56.27" />
                    <SPLIT distance="350" swimtime="00:04:38.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" points="371" reactiontime="+85" swimtime="00:03:07.31" resultid="42007" heatid="45030" lane="7" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.32" />
                    <SPLIT distance="100" swimtime="00:01:35.29" />
                    <SPLIT distance="150" swimtime="00:02:22.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="464" reactiontime="+80" swimtime="00:06:07.97" resultid="42008" heatid="45061" lane="4" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="100" swimtime="00:01:18.15" />
                    <SPLIT distance="150" swimtime="00:02:07.96" />
                    <SPLIT distance="200" swimtime="00:02:57.17" />
                    <SPLIT distance="250" swimtime="00:03:50.99" />
                    <SPLIT distance="300" swimtime="00:04:44.91" />
                    <SPLIT distance="350" swimtime="00:05:26.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Carlos" lastname="Carvalho" birthdate="1990-03-22" gender="M" nation="POR" license="25338" swrid="4074043" athleteid="42009">
              <RESULTS>
                <RESULT eventid="1058" points="402" swimtime="00:11:01.50" resultid="42010" heatid="45085" lane="8" entrytime="00:11:07.87">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.94" />
                    <SPLIT distance="200" swimtime="00:02:39.29" />
                    <SPLIT distance="300" swimtime="00:04:01.80" />
                    <SPLIT distance="400" swimtime="00:05:25.87" />
                    <SPLIT distance="500" swimtime="00:06:50.55" />
                    <SPLIT distance="600" swimtime="00:08:16.00" />
                    <SPLIT distance="700" swimtime="00:09:40.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2622" points="570" reactiontime="+88" swimtime="00:02:52.99" resultid="42011" heatid="44879" lane="7" entrytime="00:02:50.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                    <SPLIT distance="100" swimtime="00:01:22.68" />
                    <SPLIT distance="150" swimtime="00:02:08.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="554" reactiontime="+85" swimtime="00:02:40.21" resultid="42012" heatid="44982" lane="8" entrytime="00:02:37.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                    <SPLIT distance="100" swimtime="00:01:16.41" />
                    <SPLIT distance="150" swimtime="00:02:01.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="577" reactiontime="+81" swimtime="00:01:16.74" resultid="42013" heatid="44999" lane="7" entrytime="00:01:17.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" status="DNS" swimtime="00:00:00.00" resultid="42014" heatid="45062" lane="2" entrytime="00:05:40.65" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Boavida" lastname="Ferreira" birthdate="1991-06-16" gender="M" nation="POR" license="201323" swrid="5168030" athleteid="42021">
              <RESULTS>
                <RESULT eventid="2537" status="DNS" swimtime="00:00:00.00" resultid="42022" heatid="44887" lane="4" entrytime="00:01:19.00" />
                <RESULT eventid="2507" status="DNS" swimtime="00:00:00.00" resultid="42023" heatid="45094" lane="6" entrytime="00:02:30.70" />
                <RESULT eventid="2218" status="DNS" swimtime="00:00:00.00" resultid="42024" heatid="44920" lane="3" entrytime="00:02:54.20" />
                <RESULT eventid="2415" status="DNS" swimtime="00:00:00.00" resultid="42025" heatid="45112" lane="7" entrytime="00:01:05.60" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="42026" heatid="45043" lane="5" entrytime="00:00:28.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo Humberto" lastname="Viegas" birthdate="1982-09-07" gender="M" nation="POR" license="213223" swrid="5448485" athleteid="42057">
              <RESULTS>
                <RESULT eventid="2537" points="251" reactiontime="+83" swimtime="00:01:33.57" resultid="42058" heatid="44886" lane="7" entrytime="00:01:37.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="254" reactiontime="+81" swimtime="00:03:02.51" resultid="42059" heatid="45093" lane="1" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.50" />
                    <SPLIT distance="100" swimtime="00:01:21.41" />
                    <SPLIT distance="150" swimtime="00:02:10.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="304" reactiontime="+87" swimtime="00:03:17.95" resultid="42060" heatid="44919" lane="7" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.18" />
                    <SPLIT distance="100" swimtime="00:01:37.01" />
                    <SPLIT distance="150" swimtime="00:02:28.54" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="809 - Movimento alternado de pernas durante o percurso - SW 8.3" eventid="2385" reactiontime="+83" status="DSQ" swimtime="00:03:11.55" resultid="42061" heatid="44978" lane="2" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                    <SPLIT distance="100" swimtime="00:01:31.82" />
                    <SPLIT distance="150" swimtime="00:02:26.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="284" reactiontime="+80" swimtime="00:06:29.90" resultid="42062" heatid="45129" lane="2" entrytime="00:05:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.25" />
                    <SPLIT distance="100" swimtime="00:01:25.23" />
                    <SPLIT distance="150" swimtime="00:02:14.47" />
                    <SPLIT distance="200" swimtime="00:03:05.68" />
                    <SPLIT distance="250" swimtime="00:03:57.60" />
                    <SPLIT distance="300" swimtime="00:04:50.27" />
                    <SPLIT distance="350" swimtime="00:05:41.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Antonio" lastname="Pereira" birthdate="1960-03-08" gender="M" nation="POR" license="201325" swrid="5168048" athleteid="42036">
              <RESULTS>
                <RESULT eventid="2537" points="209" reactiontime="+91" swimtime="00:02:04.50" resultid="42037" heatid="44884" lane="4" entrytime="00:02:07.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="239" reactiontime="+96" swimtime="00:03:45.14" resultid="42038" heatid="45091" lane="1" entrytime="00:03:33.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.08" />
                    <SPLIT distance="100" swimtime="00:01:39.83" />
                    <SPLIT distance="150" swimtime="00:02:40.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="286" reactiontime="+90" swimtime="00:01:32.53" resultid="42039" heatid="45106" lane="8" entrytime="00:01:28.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="267" reactiontime="+81" swimtime="00:00:51.06" resultid="42040" heatid="45016" lane="1" entrytime="00:00:53.03" entrycourse="LCM" />
                <RESULT eventid="2652" points="342" reactiontime="+91" swimtime="00:00:39.06" resultid="42041" heatid="45036" lane="1" entrytime="00:00:38.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabel Xavier" lastname="Lobo" birthdate="1976-04-06" gender="F" nation="POR" license="123662" swrid="4763858" athleteid="42027">
              <RESULTS>
                <RESULT eventid="1060" points="273" swimtime="00:14:54.59" resultid="42028" heatid="45076" lane="5" entrytime="00:14:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.71" />
                    <SPLIT distance="200" swimtime="00:03:35.77" />
                    <SPLIT distance="300" swimtime="00:05:27.31" />
                    <SPLIT distance="400" swimtime="00:07:20.55" />
                    <SPLIT distance="500" swimtime="00:09:14.03" />
                    <SPLIT distance="600" swimtime="00:11:07.76" />
                    <SPLIT distance="700" swimtime="00:13:02.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2173" points="307" swimtime="00:04:13.35" resultid="42029" heatid="45087" lane="5" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.73" />
                    <SPLIT distance="100" swimtime="00:02:01.26" />
                    <SPLIT distance="150" swimtime="00:03:07.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2308" points="235" reactiontime="+101" swimtime="00:04:17.80" resultid="42030" heatid="44913" lane="5" entrytime="00:04:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.52" />
                    <SPLIT distance="100" swimtime="00:02:03.69" />
                    <SPLIT distance="150" swimtime="00:03:11.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="287" reactiontime="+95" swimtime="00:07:11.07" resultid="42031" heatid="45010" lane="2" entrytime="00:07:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.18" />
                    <SPLIT distance="100" swimtime="00:01:39.01" />
                    <SPLIT distance="150" swimtime="00:02:33.51" />
                    <SPLIT distance="200" swimtime="00:03:28.66" />
                    <SPLIT distance="250" swimtime="00:04:24.18" />
                    <SPLIT distance="300" swimtime="00:05:19.83" />
                    <SPLIT distance="350" swimtime="00:06:16.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Filipe" lastname="Almeida" birthdate="1966-07-27" gender="M" nation="POR" license="201324" swrid="5168018" athleteid="41998">
              <RESULTS>
                <RESULT eventid="2218" points="246" reactiontime="+118" swimtime="00:04:00.97" resultid="41999" heatid="44918" lane="8" entrytime="00:03:50.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.72" />
                    <SPLIT distance="100" swimtime="00:01:57.89" />
                    <SPLIT distance="150" swimtime="00:02:59.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="320" reactiontime="+103" swimtime="00:00:45.37" resultid="42000" heatid="44944" lane="5" entrytime="00:00:43.81" />
                <RESULT eventid="2385" points="328" reactiontime="+97" swimtime="00:03:42.04" resultid="42001" heatid="44977" lane="8" entrytime="00:03:39.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.73" />
                    <SPLIT distance="100" swimtime="00:01:52.65" />
                    <SPLIT distance="150" swimtime="00:02:51.71" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="403 - Falsa partida - SW 4.4" eventid="2567" reactiontime="+86" status="DSQ" swimtime="00:04:29.06" resultid="42002" heatid="45028" lane="4" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.89" />
                    <SPLIT distance="100" swimtime="00:02:11.11" />
                    <SPLIT distance="150" swimtime="00:03:20.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="328" reactiontime="+101" swimtime="00:07:59.95" resultid="42003" heatid="45059" lane="3" entrytime="00:07:56.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.48" />
                    <SPLIT distance="100" swimtime="00:01:59.82" />
                    <SPLIT distance="150" swimtime="00:03:04.43" />
                    <SPLIT distance="200" swimtime="00:04:07.41" />
                    <SPLIT distance="250" swimtime="00:05:13.73" />
                    <SPLIT distance="300" swimtime="00:06:15.32" />
                    <SPLIT distance="350" swimtime="00:07:08.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Filipe" lastname="Pinto" birthdate="1982-09-13" gender="M" nation="POR" license="207564" swrid="4532500" athleteid="42048">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="42049" heatid="45085" lane="1" entrytime="00:11:07.00" />
                <RESULT eventid="2385" points="612" reactiontime="+73" swimtime="00:02:35.57" resultid="42050" heatid="44981" lane="5" entrytime="00:02:38.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                    <SPLIT distance="100" swimtime="00:01:11.16" />
                    <SPLIT distance="150" swimtime="00:01:55.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="598" reactiontime="+74" swimtime="00:05:38.18" resultid="42051" heatid="45062" lane="1" entrytime="00:05:42.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:11.07" />
                    <SPLIT distance="150" swimtime="00:01:55.47" />
                    <SPLIT distance="200" swimtime="00:02:38.42" />
                    <SPLIT distance="250" swimtime="00:03:26.66" />
                    <SPLIT distance="300" swimtime="00:04:16.16" />
                    <SPLIT distance="350" swimtime="00:04:57.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCB" nation="POR" region="ANMIN" clubid="42998" swrid="65807" name="Sporting Clube de Braga" shortname="Braga">
          <ATHLETES>
            <ATHLETE firstname="Nuno Carlos" lastname="Albuquerque" birthdate="1964-07-19" gender="M" nation="POR" license="210412" swrid="5361434" athleteid="43068">
              <RESULTS>
                <RESULT eventid="1058" points="271" swimtime="00:14:35.34" resultid="43069" heatid="45081" lane="1" entrytime="00:15:31.31">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.00" />
                    <SPLIT distance="200" swimtime="00:03:29.86" />
                    <SPLIT distance="300" swimtime="00:05:21.08" />
                    <SPLIT distance="400" swimtime="00:07:12.34" />
                    <SPLIT distance="500" swimtime="00:09:04.42" />
                    <SPLIT distance="600" swimtime="00:10:55.39" />
                    <SPLIT distance="700" swimtime="00:12:46.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="236" reactiontime="+109" swimtime="00:00:45.73" resultid="43070" heatid="44893" lane="5" entrytime="00:00:48.51" entrycourse="SCM" />
                <RESULT eventid="2323" points="194" reactiontime="+88" swimtime="00:01:51.57" resultid="43071" heatid="44925" lane="5" entrytime="00:02:02.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="269" reactiontime="+101" swimtime="00:07:07.72" resultid="43072" heatid="45126" lane="8" entrytime="00:07:39.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.45" />
                    <SPLIT distance="100" swimtime="00:01:37.84" />
                    <SPLIT distance="150" swimtime="00:02:31.36" />
                    <SPLIT distance="200" swimtime="00:03:27.15" />
                    <SPLIT distance="250" swimtime="00:04:21.38" />
                    <SPLIT distance="300" swimtime="00:05:17.74" />
                    <SPLIT distance="350" swimtime="00:06:12.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="283" reactiontime="+83" swimtime="00:00:40.53" resultid="43073" heatid="45035" lane="8" entrytime="00:00:42.20" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago Nuno" lastname="Pimentel" birthdate="1985-08-02" gender="M" nation="POR" license="212448" swrid="5429852" athleteid="43088">
              <RESULTS>
                <RESULT comment="403 - Falsa partida - SW 4.4" eventid="2188" reactiontime="+88" status="DSQ" swimtime="00:00:45.31" resultid="43089" heatid="44945" lane="3" entrytime="00:00:42.00" entrycourse="SCM" />
                <RESULT eventid="2445" points="279" reactiontime="+91" swimtime="00:01:41.63" resultid="43090" heatid="44995" lane="8" entrytime="00:01:40.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="247" reactiontime="+96" swimtime="00:06:48.63" resultid="43091" heatid="45126" lane="4" entrytime="00:06:58.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.64" />
                    <SPLIT distance="100" swimtime="00:01:29.76" />
                    <SPLIT distance="150" swimtime="00:02:20.29" />
                    <SPLIT distance="200" swimtime="00:03:13.22" />
                    <SPLIT distance="250" swimtime="00:04:07.84" />
                    <SPLIT distance="300" swimtime="00:05:02.54" />
                    <SPLIT distance="350" swimtime="00:05:57.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="237" reactiontime="+97" swimtime="00:07:39.86" resultid="43092" heatid="45060" lane="4" entrytime="00:06:31.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.12" />
                    <SPLIT distance="100" swimtime="00:01:44.80" />
                    <SPLIT distance="150" swimtime="00:02:46.87" />
                    <SPLIT distance="200" swimtime="00:03:49.67" />
                    <SPLIT distance="250" swimtime="00:04:51.68" />
                    <SPLIT distance="300" swimtime="00:05:53.37" />
                    <SPLIT distance="350" swimtime="00:06:47.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gilberto Luis" lastname="Ferreira" birthdate="1985-02-07" gender="M" nation="POR" license="211915" swrid="5425454" athleteid="43074">
              <RESULTS>
                <RESULT eventid="2507" points="301" reactiontime="+94" swimtime="00:02:52.59" resultid="43075" heatid="45093" lane="4" entrytime="00:02:40.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                    <SPLIT distance="100" swimtime="00:01:19.65" />
                    <SPLIT distance="150" swimtime="00:02:06.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="270" reactiontime="+99" swimtime="00:03:24.19" resultid="43076" heatid="44980" lane="6" entrytime="00:02:51.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                    <SPLIT distance="100" swimtime="00:01:38.02" />
                    <SPLIT distance="150" swimtime="00:02:36.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="318" reactiontime="+89" swimtime="00:06:15.62" resultid="43077" heatid="45127" lane="3" entrytime="00:06:35.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                    <SPLIT distance="100" swimtime="00:01:28.62" />
                    <SPLIT distance="150" swimtime="00:02:17.18" />
                    <SPLIT distance="200" swimtime="00:03:06.22" />
                    <SPLIT distance="250" swimtime="00:03:54.96" />
                    <SPLIT distance="300" swimtime="00:04:43.82" />
                    <SPLIT distance="350" swimtime="00:05:32.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joana Marques" lastname="Maia" birthdate="1991-03-16" gender="F" nation="POR" license="25067" swrid="4269239" athleteid="43078">
              <RESULTS>
                <RESULT comment="Rec Nac Esc B" eventid="2173" points="873" swimtime="00:02:46.69" resultid="43079" heatid="45089" lane="5" entrytime="00:02:47.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                    <SPLIT distance="100" swimtime="00:01:18.80" />
                    <SPLIT distance="150" swimtime="00:02:02.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="715" reactiontime="+81" swimtime="00:00:36.03" resultid="43080" heatid="45103" lane="4" entrytime="00:00:36.07" entrycourse="LCM" />
                <RESULT eventid="2460" points="827" reactiontime="+79" swimtime="00:01:16.68" resultid="43081" heatid="45123" lane="4" entrytime="00:01:17.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Goncalo Goncalves" lastname="Meneses" birthdate="1992-06-06" gender="M" nation="POR" license="204349" swrid="4269434" athleteid="43082">
              <RESULTS>
                <RESULT eventid="2622" points="427" reactiontime="+95" swimtime="00:03:12.02" resultid="43083" heatid="44879" lane="6" entrytime="00:02:46.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                    <SPLIT distance="100" swimtime="00:01:29.34" />
                    <SPLIT distance="150" swimtime="00:02:20.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="417" reactiontime="+88" swimtime="00:00:38.63" resultid="43084" heatid="44949" lane="5" entrytime="00:00:35.10" entrycourse="SCM" />
                <RESULT eventid="2385" points="483" reactiontime="+90" swimtime="00:02:40.47" resultid="43085" heatid="44982" lane="3" entrytime="00:02:28.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:14.63" />
                    <SPLIT distance="150" swimtime="00:02:02.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="341" reactiontime="+97" swimtime="00:01:31.50" resultid="43086" heatid="44999" lane="1" entrytime="00:01:18.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="490" reactiontime="+91" swimtime="00:06:01.91" resultid="43087" heatid="45062" lane="3" entrytime="00:05:20.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                    <SPLIT distance="100" swimtime="00:01:15.80" />
                    <SPLIT distance="150" swimtime="00:02:04.09" />
                    <SPLIT distance="200" swimtime="00:02:50.85" />
                    <SPLIT distance="250" swimtime="00:03:43.94" />
                    <SPLIT distance="300" swimtime="00:04:38.76" />
                    <SPLIT distance="350" swimtime="00:05:20.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SFUS" nation="POR" region="ANDS" clubid="41721" swrid="68066" name="Sociedade Filarmonica Uniao Samorense" shortname="Uniao Samorense">
          <ATHLETES>
            <ATHLETE firstname="Vanessa Braga" lastname="Salvador" birthdate="1991-10-25" gender="F" nation="POR" license="11370" swrid="4074005" athleteid="41722">
              <RESULTS>
                <RESULT eventid="2338" points="713" reactiontime="+84" swimtime="00:00:32.01" resultid="41723" heatid="44892" lane="3" entrytime="00:00:31.82" entrycourse="LCM" />
                <RESULT eventid="2552" points="784" reactiontime="+83" swimtime="00:01:09.99" resultid="41724" heatid="44924" lane="6" entrytime="00:01:09.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2667" points="750" reactiontime="+92" swimtime="00:02:37.98" resultid="41725" heatid="45031" lane="4" entrytime="00:02:39.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                    <SPLIT distance="100" swimtime="00:01:13.88" />
                    <SPLIT distance="150" swimtime="00:01:54.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CAP" nation="POR" region="ANNP" clubid="41797" swrid="89149" name="Clube Aquatico Pacense" shortname="Aquatico Pacense">
          <ATHLETES>
            <ATHLETE firstname="Antonio Rafael" lastname="Bessa" birthdate="1994-03-25" gender="M" nation="POR" license="102089" swrid="4574455" athleteid="41798">
              <RESULTS>
                <RESULT eventid="2567" points="885" reactiontime="+71" swimtime="00:02:13.50" resultid="41799" heatid="45030" lane="5" entrytime="00:02:07.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.25" />
                    <SPLIT distance="100" swimtime="00:01:03.09" />
                    <SPLIT distance="150" swimtime="00:01:37.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CNMAL" nation="POR" region="ANL" clubid="41551" swrid="73262" name="Clube Natacao Masters de Almada" shortname="Masters de Almada">
          <ATHLETES>
            <ATHLETE firstname="Fernanda Maria" lastname="Santinha" birthdate="1972-05-23" gender="F" nation="POR" license="100478" swrid="4345983" athleteid="43766">
              <RESULTS>
                <RESULT eventid="1060" status="DNS" swimtime="00:00:00.00" resultid="43767" heatid="45076" lane="6" entrytime="00:14:38.30" />
                <RESULT eventid="2173" status="DNS" swimtime="00:00:00.00" resultid="43768" heatid="45087" lane="4" entrytime="00:04:08.34" />
                <RESULT eventid="2492" status="DNS" swimtime="00:00:00.00" resultid="43769" heatid="45010" lane="3" entrytime="00:07:11.12" />
                <RESULT eventid="2667" status="DNS" swimtime="00:00:00.00" resultid="43770" heatid="45031" lane="7" entrytime="00:04:21.03" />
                <RESULT eventid="2400" status="DNS" swimtime="00:00:00.00" resultid="43771" heatid="45063" lane="3" entrytime="00:08:34.91" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Henriques" lastname="Pato" birthdate="1983-08-16" gender="F" nation="POR" license="204148" swrid="5133139" athleteid="43777">
              <RESULTS>
                <RESULT eventid="2203" points="362" reactiontime="+75" swimtime="00:01:37.73" resultid="43778" heatid="44882" lane="3" entrytime="00:01:32.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="329" reactiontime="+89" swimtime="00:00:47.31" resultid="43779" heatid="45101" lane="2" entrytime="00:00:46.24" />
                <RESULT eventid="2522" points="423" reactiontime="+94" swimtime="00:00:42.68" resultid="43780" heatid="45026" lane="1" entrytime="00:00:41.33" />
                <RESULT eventid="2430" points="468" reactiontime="+84" swimtime="00:00:34.55" resultid="43781" heatid="45070" lane="4" entrytime="00:00:34.31" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Goncalves" lastname="Vasconcelos" birthdate="1964-12-19" gender="F" nation="POR" license="130670" swrid="5003489" athleteid="43755">
              <RESULTS>
                <RESULT eventid="2338" points="234" reactiontime="+110" swimtime="00:00:51.62" resultid="43756" heatid="44890" lane="7" entrytime="00:00:50.87" />
                <RESULT eventid="2552" points="203" reactiontime="+114" swimtime="00:02:04.33" resultid="43757" heatid="44922" lane="4" entrytime="00:02:06.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="301" reactiontime="+120" swimtime="00:01:34.93" resultid="43758" heatid="44954" lane="1" entrytime="00:01:36.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="345" reactiontime="+115" swimtime="00:00:42.20" resultid="43759" heatid="45068" lane="1" entrytime="00:00:42.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Dinis" lastname="Freitas" birthdate="1983-10-28" gender="M" nation="POR" license="204149" swrid="5133138" athleteid="43788">
              <RESULTS>
                <RESULT eventid="1058" points="244" swimtime="00:14:16.97" resultid="43789" heatid="45081" lane="5" entrytime="00:14:03.34">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.29" />
                    <SPLIT distance="200" swimtime="00:03:22.04" />
                    <SPLIT distance="300" swimtime="00:05:12.34" />
                    <SPLIT distance="400" swimtime="00:07:06.17" />
                    <SPLIT distance="500" swimtime="00:08:58.97" />
                    <SPLIT distance="600" swimtime="00:10:52.02" />
                    <SPLIT distance="700" swimtime="00:12:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2622" points="282" reactiontime="+90" swimtime="00:03:50.62" resultid="43790" heatid="44876" lane="1" entrytime="00:03:33.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.53" />
                    <SPLIT distance="100" swimtime="00:01:52.82" />
                    <SPLIT distance="150" swimtime="00:02:54.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="228" reactiontime="+87" swimtime="00:00:41.76" resultid="43791" heatid="44894" lane="7" entrytime="00:00:45.41" />
                <RESULT eventid="2218" points="181" reactiontime="+91" swimtime="00:03:55.36" resultid="43792" heatid="44918" lane="3" entrytime="00:03:37.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.17" />
                    <SPLIT distance="100" swimtime="00:01:54.32" />
                    <SPLIT distance="150" swimtime="00:02:56.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="275" reactiontime="+91" swimtime="00:00:44.91" resultid="43793" heatid="44944" lane="3" entrytime="00:00:43.85" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos Augusto" lastname="Correia" birthdate="1952-03-18" gender="M" nation="POR" license="100466" swrid="4345463" athleteid="43127">
              <RESULTS>
                <RESULT eventid="1058" points="403" swimtime="00:14:35.43" resultid="43128" heatid="45080" lane="4" entrytime="00:14:00.98">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.77" />
                    <SPLIT distance="200" swimtime="00:03:38.39" />
                    <SPLIT distance="300" swimtime="00:05:29.60" />
                    <SPLIT distance="400" swimtime="00:07:20.73" />
                    <SPLIT distance="500" swimtime="00:09:11.46" />
                    <SPLIT distance="600" swimtime="00:11:02.31" />
                    <SPLIT distance="700" swimtime="00:12:51.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2537" points="215" reactiontime="+85" swimtime="00:02:03.07" resultid="43129" heatid="44885" lane="1" entrytime="00:02:01.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="387" reactiontime="+118" swimtime="00:03:20.91" resultid="43130" heatid="45092" lane="8" entrytime="00:03:13.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                    <SPLIT distance="100" swimtime="00:01:35.61" />
                    <SPLIT distance="150" swimtime="00:02:29.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="304" reactiontime="+111" swimtime="00:04:06.12" resultid="43131" heatid="44976" lane="7" entrytime="00:03:57.08">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.21" />
                    <SPLIT distance="100" swimtime="00:02:05.18" />
                    <SPLIT distance="150" swimtime="00:03:16.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="419" reactiontime="+116" swimtime="00:06:59.82" resultid="43132" heatid="45127" lane="1" entrytime="00:06:44.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.86" />
                    <SPLIT distance="100" swimtime="00:01:39.91" />
                    <SPLIT distance="150" swimtime="00:02:33.57" />
                    <SPLIT distance="200" swimtime="00:03:29.01" />
                    <SPLIT distance="250" swimtime="00:04:21.50" />
                    <SPLIT distance="300" swimtime="00:05:15.88" />
                    <SPLIT distance="350" swimtime="00:06:07.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Gabriel" lastname="David" birthdate="1987-08-12" gender="M" nation="BRA" license="210595" swrid="5145168" athleteid="43782">
              <RESULTS>
                <RESULT eventid="2682" points="410" reactiontime="+72" swimtime="00:00:33.67" resultid="43783" heatid="44897" lane="2" entrytime="00:00:34.25" />
                <RESULT eventid="2188" points="397" reactiontime="+80" swimtime="00:00:39.16" resultid="43784" heatid="44946" lane="4" entrytime="00:00:39.65" />
                <RESULT eventid="2415" points="399" reactiontime="+79" swimtime="00:01:09.01" resultid="43785" heatid="45111" lane="3" entrytime="00:01:07.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="373" reactiontime="+77" swimtime="00:01:28.75" resultid="43786" heatid="44997" lane="2" entrytime="00:01:28.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="467" reactiontime="+76" swimtime="00:00:29.96" resultid="43787" heatid="45042" lane="5" entrytime="00:00:29.76" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Manuel" lastname="Santinha" birthdate="1969-12-31" gender="M" nation="POR" license="100477" swrid="4345982" athleteid="43760">
              <RESULTS>
                <RESULT eventid="1058" points="270" swimtime="00:14:11.93" resultid="43761" heatid="45082" lane="1" entrytime="00:13:48.78">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.55" />
                    <SPLIT distance="200" swimtime="00:03:31.36" />
                    <SPLIT distance="300" swimtime="00:05:19.51" />
                    <SPLIT distance="400" swimtime="00:07:08.53" />
                    <SPLIT distance="500" swimtime="00:08:56.74" />
                    <SPLIT distance="600" swimtime="00:10:43.26" />
                    <SPLIT distance="700" swimtime="00:12:29.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2622" points="333" reactiontime="+110" swimtime="00:03:50.73" resultid="43762" heatid="44875" lane="7" entrytime="00:03:44.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.65" />
                    <SPLIT distance="100" swimtime="00:01:56.94" />
                    <SPLIT distance="150" swimtime="00:02:57.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="341" reactiontime="+98" swimtime="00:00:44.54" resultid="43763" heatid="44944" lane="6" entrytime="00:00:44.08" />
                <RESULT eventid="2263" points="272" reactiontime="+110" swimtime="00:06:52.23" resultid="43764" heatid="45127" lane="8" entrytime="00:06:50.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.66" />
                    <SPLIT distance="100" swimtime="00:01:38.24" />
                    <SPLIT distance="150" swimtime="00:02:31.12" />
                    <SPLIT distance="200" swimtime="00:03:23.85" />
                    <SPLIT distance="250" swimtime="00:04:17.22" />
                    <SPLIT distance="300" swimtime="00:05:09.43" />
                    <SPLIT distance="350" swimtime="00:06:02.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="361" reactiontime="+93" swimtime="00:01:41.78" resultid="43765" heatid="44994" lane="4" entrytime="00:01:40.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina Isabel" lastname="Mendes" birthdate="1968-08-22" gender="F" nation="POR" license="106063" swrid="4345754" athleteid="43750">
              <RESULTS>
                <RESULT eventid="2552" points="178" reactiontime="+99" swimtime="00:02:06.91" resultid="43751" heatid="44923" lane="8" entrytime="00:02:03.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="367" reactiontime="+105" swimtime="00:00:51.25" resultid="43752" heatid="45100" lane="2" entrytime="00:00:49.92" />
                <RESULT eventid="2460" points="380" reactiontime="+107" swimtime="00:01:54.55" resultid="43753" heatid="45119" lane="6" entrytime="00:02:00.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="338" reactiontime="+96" swimtime="00:00:40.77" resultid="43754" heatid="45069" lane="8" entrytime="00:00:39.14" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo Felipi" lastname="Costa" birthdate="1979-11-27" gender="M" nation="BRA" license="213752" swrid="5455231" athleteid="43794">
              <RESULTS>
                <RESULT eventid="2415" points="457" reactiontime="+90" swimtime="00:01:10.51" resultid="43795" heatid="45109" lane="6" entrytime="00:01:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="402" reactiontime="+72" swimtime="00:00:38.48" resultid="43796" heatid="45018" lane="7" entrytime="00:00:43.00" />
                <RESULT eventid="2652" points="569" reactiontime="+93" swimtime="00:00:29.66" resultid="43797" heatid="45041" lane="2" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos Jorge" lastname="Oliveira" birthdate="1964-02-16" gender="M" nation="POR" license="11360" swrid="4800238" athleteid="43798">
              <RESULTS>
                <RESULT eventid="1058" points="529" swimtime="00:11:41.13" resultid="43799" heatid="45084" lane="5" entrytime="00:11:16.51">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.91" />
                    <SPLIT distance="200" swimtime="00:02:48.72" />
                    <SPLIT distance="300" swimtime="00:04:18.38" />
                    <SPLIT distance="400" swimtime="00:05:47.58" />
                    <SPLIT distance="500" swimtime="00:07:16.50" />
                    <SPLIT distance="600" swimtime="00:08:45.14" />
                    <SPLIT distance="700" swimtime="00:10:13.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2537" points="528" reactiontime="+67" swimtime="00:01:24.44" resultid="43800" heatid="44887" lane="2" entrytime="00:01:27.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="500" reactiontime="+107" swimtime="00:00:35.64" resultid="43801" heatid="44896" lane="3" entrytime="00:00:36.16" />
                <RESULT eventid="2218" points="533" reactiontime="+74" swimtime="00:03:06.16" resultid="43802" heatid="44920" lane="1" entrytime="00:03:05.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.39" />
                    <SPLIT distance="100" swimtime="00:01:29.13" />
                    <SPLIT distance="150" swimtime="00:02:18.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2323" points="322" reactiontime="+100" swimtime="00:01:34.20" resultid="43803" heatid="44926" lane="6" entrytime="00:01:38.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joana Pereira" lastname="Barbara" birthdate="1987-01-06" gender="F" nation="POR" license="13948" swrid="4062691" athleteid="43772">
              <RESULTS>
                <RESULT eventid="2607" points="610" reactiontime="+83" swimtime="00:00:37.99" resultid="43773" heatid="45103" lane="3" entrytime="00:00:36.74" />
                <RESULT eventid="2637" points="565" reactiontime="+82" swimtime="00:01:10.46" resultid="43774" heatid="44957" lane="2" entrytime="00:01:08.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="506" reactiontime="+86" swimtime="00:01:30.31" resultid="43775" heatid="45123" lane="3" entrytime="00:01:25.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="559" reactiontime="+78" swimtime="00:00:32.12" resultid="43776" heatid="45073" lane="8" entrytime="00:00:30.37" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carla Filomena" lastname="Peixe" birthdate="1963-06-19" gender="F" nation="POR" license="14184" swrid="4575460" athleteid="43746">
              <RESULTS>
                <RESULT eventid="2607" points="367" reactiontime="+112" swimtime="00:00:52.75" resultid="43747" heatid="45099" lane="1" entrytime="00:00:52.58" />
                <RESULT eventid="2460" points="373" reactiontime="+106" swimtime="00:01:57.75" resultid="43748" heatid="45120" lane="3" entrytime="00:01:50.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="398" reactiontime="+99" swimtime="00:00:40.24" resultid="43749" heatid="45068" lane="6" entrytime="00:00:39.80" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Madalena" lastname="Caninas" birthdate="1963-11-20" gender="F" nation="POR" license="108658" swrid="4345423" athleteid="43121">
              <RESULTS>
                <RESULT eventid="1060" points="232" swimtime="00:16:24.31" resultid="43122" heatid="45076" lane="2" entrytime="00:15:11.36">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:51.22" />
                    <SPLIT distance="200" swimtime="00:03:56.29" />
                    <SPLIT distance="300" swimtime="00:06:02.97" />
                    <SPLIT distance="400" swimtime="00:08:10.73" />
                    <SPLIT distance="500" swimtime="00:10:16.98" />
                    <SPLIT distance="600" swimtime="00:12:22.30" />
                    <SPLIT distance="700" swimtime="00:14:25.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2338" points="164" reactiontime="+116" swimtime="00:00:58.09" resultid="43123" heatid="44889" lane="3" entrytime="00:01:00.20" />
                <RESULT eventid="2278" points="324" reactiontime="+107" swimtime="00:03:23.39" resultid="43124" heatid="44903" lane="8" entrytime="00:03:28.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.90" />
                    <SPLIT distance="100" swimtime="00:01:37.26" />
                    <SPLIT distance="150" swimtime="00:02:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="215" reactiontime="+119" swimtime="00:04:25.21" resultid="43125" heatid="44971" lane="3" entrytime="00:04:27.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.25" />
                    <SPLIT distance="100" swimtime="00:02:14.62" />
                    <SPLIT distance="150" swimtime="00:03:32.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="269" reactiontime="+113" swimtime="00:07:30.25" resultid="43126" heatid="45010" lane="1" entrytime="00:07:25.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.84" />
                    <SPLIT distance="100" swimtime="00:01:43.55" />
                    <SPLIT distance="150" swimtime="00:02:42.78" />
                    <SPLIT distance="200" swimtime="00:03:43.88" />
                    <SPLIT distance="250" swimtime="00:04:43.28" />
                    <SPLIT distance="300" swimtime="00:05:43.39" />
                    <SPLIT distance="350" swimtime="00:06:40.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jorge Manuel" lastname="Roque" birthdate="1990-05-14" gender="M" nation="POR" license="10760" swrid="4074217" athleteid="43740">
              <RESULTS>
                <RESULT eventid="2682" points="808" reactiontime="+74" swimtime="00:00:26.86" resultid="43741" heatid="44901" lane="4" entrytime="00:00:26.56" />
                <RESULT eventid="2507" points="685" reactiontime="+79" swimtime="00:02:11.23" resultid="43742" heatid="45096" lane="4" entrytime="00:02:04.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.17" />
                    <SPLIT distance="100" swimtime="00:01:03.82" />
                    <SPLIT distance="150" swimtime="00:01:38.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2323" points="796" reactiontime="+80" swimtime="00:01:01.16" resultid="43743" heatid="44930" lane="4" entrytime="00:00:58.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="659" reactiontime="+74" swimtime="00:00:58.42" resultid="43744" heatid="45116" lane="6" entrytime="00:00:55.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="720" reactiontime="+79" swimtime="00:00:25.94" resultid="43745" heatid="45048" lane="3" entrytime="00:00:25.45" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCE" nation="POR" region="ANCNP" clubid="42741" swrid="65808" name="Sporting Clube de Espinho" shortname="Sporting de Espinho">
          <ATHLETES>
            <ATHLETE firstname="Fabio" lastname="Floriano" birthdate="1963-10-07" gender="M" nation="POR" license="207665" swrid="5297527" athleteid="42754">
              <RESULTS>
                <RESULT eventid="2188" status="DNS" swimtime="00:00:00.00" resultid="42755" heatid="44945" lane="8" entrytime="00:00:43.19" entrycourse="LCM" />
                <RESULT eventid="2445" status="DNS" swimtime="00:00:00.00" resultid="42756" heatid="44995" lane="1" entrytime="00:01:40.44" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Monteiro" lastname="Canelas" birthdate="1950-01-26" gender="M" nation="POR" license="148547" swrid="5100108" athleteid="42742">
              <RESULTS>
                <RESULT eventid="2682" points="260" reactiontime="+97" swimtime="00:00:49.47" resultid="42743" heatid="44894" lane="8" entrytime="00:00:46.55" entrycourse="LCM" />
                <RESULT eventid="2323" points="246" reactiontime="+112" swimtime="00:02:04.51" resultid="42744" heatid="44926" lane="1" entrytime="00:01:53.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="294" reactiontime="+112" swimtime="00:04:30.56" resultid="42745" heatid="44975" lane="5" entrytime="00:04:09.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.99" />
                    <SPLIT distance="100" swimtime="00:02:19.00" />
                    <SPLIT distance="150" swimtime="00:03:28.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="173" reactiontime="+112" swimtime="00:01:02.61" resultid="42746" heatid="45015" lane="8" entrytime="00:01:01.47" entrycourse="LCM" />
                <RESULT eventid="2248" points="292" reactiontime="+114" swimtime="00:10:03.29" resultid="42747" heatid="45058" lane="5" entrytime="00:09:23.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.38" />
                    <SPLIT distance="100" swimtime="00:02:13.57" />
                    <SPLIT distance="150" swimtime="00:03:55.59" />
                    <SPLIT distance="200" swimtime="00:05:23.45" />
                    <SPLIT distance="250" swimtime="00:06:35.73" />
                    <SPLIT distance="300" swimtime="00:07:51.20" />
                    <SPLIT distance="350" swimtime="00:09:00.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Domingos Jose" lastname="Ferreira" birthdate="1954-11-05" gender="M" nation="POR" license="209351" swrid="5336707" athleteid="42748">
              <RESULTS>
                <RESULT eventid="2507" points="370" reactiontime="+104" swimtime="00:03:23.90" resultid="42749" heatid="45091" lane="4" entrytime="00:03:18.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:01:32.10" />
                    <SPLIT distance="150" swimtime="00:02:28.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="284" reactiontime="+110" swimtime="00:00:52.45" resultid="42750" heatid="44940" lane="7" entrytime="00:00:51.04" entrycourse="LCM" />
                <RESULT eventid="2415" points="305" reactiontime="+114" swimtime="00:01:33.24" resultid="42751" heatid="45106" lane="2" entrytime="00:01:27.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="383" reactiontime="+109" swimtime="00:07:12.73" resultid="42752" heatid="45126" lane="6" entrytime="00:07:04.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                    <SPLIT distance="100" swimtime="00:01:37.98" />
                    <SPLIT distance="150" swimtime="00:02:34.98" />
                    <SPLIT distance="200" swimtime="00:03:30.66" />
                    <SPLIT distance="250" swimtime="00:04:27.88" />
                    <SPLIT distance="300" swimtime="00:05:24.44" />
                    <SPLIT distance="350" swimtime="00:06:20.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="318" reactiontime="+109" swimtime="00:00:41.55" resultid="42753" heatid="45035" lane="5" entrytime="00:00:39.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Manuela" lastname="Oliveira" birthdate="1974-11-07" gender="F" nation="POR" license="208451" swrid="5326883" athleteid="42757">
              <RESULTS>
                <RESULT eventid="2607" points="356" reactiontime="+68" swimtime="00:00:51.05" resultid="42758" heatid="45100" lane="7" entrytime="00:00:49.95" entrycourse="LCM" />
                <RESULT eventid="2637" points="324" reactiontime="+81" swimtime="00:01:27.21" resultid="42759" heatid="44954" lane="3" entrytime="00:01:31.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="333" swimtime="00:01:55.54" resultid="42760" heatid="45120" lane="2" entrytime="00:01:52.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="FCP" nation="POR" region="ANNP" clubid="41930" swrid="78213" name="Futebol Clube do Porto" shortname="Porto">
          <ATHLETES>
            <ATHLETE firstname="Joao Filipe" lastname="Carvalho" birthdate="1987-07-29" gender="M" nation="POR" license="23026" swrid="4064518" athleteid="42104">
              <RESULTS>
                <RESULT eventid="2415" points="745" reactiontime="+70" swimtime="00:00:56.07" resultid="42105" heatid="45116" lane="4" entrytime="00:00:49.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="583" reactiontime="+80" swimtime="00:00:31.14" resultid="42106" heatid="45022" lane="7" entrytime="00:00:32.25" />
                <RESULT eventid="2652" points="767" reactiontime="+71" swimtime="00:00:25.39" resultid="42107" heatid="45048" lane="5" entrytime="00:00:25.28" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Manuel" lastname="Friaes" birthdate="1965-01-13" gender="F" nation="POR" license="204549" swrid="5207367" athleteid="42131">
              <RESULTS>
                <RESULT eventid="2203" points="487" reactiontime="+79" swimtime="00:01:39.30" resultid="42132" heatid="44881" lane="6" entrytime="00:01:52.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2338" points="533" reactiontime="+90" swimtime="00:00:39.25" resultid="42133" heatid="44890" lane="5" entrytime="00:00:42.61" entrycourse="LCM" />
                <RESULT eventid="2308" points="439" reactiontime="+96" swimtime="00:03:39.66" resultid="42134" heatid="44913" lane="3" entrytime="00:04:13.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.90" />
                    <SPLIT distance="100" swimtime="00:01:50.25" />
                    <SPLIT distance="150" swimtime="00:02:46.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2552" points="361" reactiontime="+104" swimtime="00:01:42.70" resultid="42135" heatid="44923" lane="2" entrytime="00:01:59.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2667" points="335" reactiontime="+105" swimtime="00:03:56.26" resultid="42136" heatid="45031" lane="1" entrytime="00:04:38.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.57" />
                    <SPLIT distance="100" swimtime="00:01:52.92" />
                    <SPLIT distance="150" swimtime="00:02:56.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mario Jorge" lastname="Barros" birthdate="1956-06-06" gender="M" nation="POR" license="128252" swrid="4913068" athleteid="42098">
              <RESULTS>
                <RESULT eventid="2622" points="573" reactiontime="+94" swimtime="00:03:45.73" resultid="42099" heatid="44875" lane="5" entrytime="00:03:40.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.34" />
                    <SPLIT distance="100" swimtime="00:01:52.54" />
                    <SPLIT distance="150" swimtime="00:02:52.10" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="403 - Falsa partida - SW 4.4" eventid="2218" reactiontime="+85" status="DSQ" swimtime="00:03:52.44" resultid="42100" heatid="44918" lane="7" entrytime="00:03:47.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.35" />
                    <SPLIT distance="100" swimtime="00:01:56.03" />
                    <SPLIT distance="150" swimtime="00:02:57.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="458" reactiontime="+96" swimtime="00:00:44.77" resultid="42101" heatid="44943" lane="6" entrytime="00:00:44.96" entrycourse="LCM" />
                <RESULT eventid="2385" points="406" reactiontime="+102" swimtime="00:03:43.52" resultid="42102" heatid="44976" lane="2" entrytime="00:03:48.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.15" />
                    <SPLIT distance="100" swimtime="00:01:54.88" />
                    <SPLIT distance="150" swimtime="00:02:53.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="419" reactiontime="+105" swimtime="00:08:24.01" resultid="42103" heatid="45059" lane="2" entrytime="00:08:11.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.17" />
                    <SPLIT distance="100" swimtime="00:02:03.14" />
                    <SPLIT distance="150" swimtime="00:03:11.62" />
                    <SPLIT distance="200" swimtime="00:04:16.75" />
                    <SPLIT distance="250" swimtime="00:05:23.10" />
                    <SPLIT distance="300" swimtime="00:06:26.80" />
                    <SPLIT distance="350" swimtime="00:07:27.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gisela Barbosa" lastname="Coutinho" birthdate="1975-01-18" gender="F" nation="POR" license="211764" swrid="5418285" athleteid="42119">
              <RESULTS>
                <RESULT eventid="2308" points="734" reactiontime="+82" swimtime="00:02:56.39" resultid="42120" heatid="44915" lane="4" entrytime="00:02:25.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:22.77" />
                    <SPLIT distance="150" swimtime="00:02:09.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="670" reactiontime="+101" swimtime="00:02:53.65" resultid="42121" heatid="44972" lane="3" entrytime="00:03:25.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                    <SPLIT distance="100" swimtime="00:01:19.49" />
                    <SPLIT distance="150" swimtime="00:02:11.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="638" reactiontime="+106" swimtime="00:05:30.17" resultid="42122" heatid="45012" lane="1" entrytime="00:06:25.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                    <SPLIT distance="100" swimtime="00:01:17.84" />
                    <SPLIT distance="150" swimtime="00:01:59.36" />
                    <SPLIT distance="200" swimtime="00:02:42.03" />
                    <SPLIT distance="250" swimtime="00:03:24.26" />
                    <SPLIT distance="300" swimtime="00:04:07.69" />
                    <SPLIT distance="350" swimtime="00:04:49.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="576" reactiontime="+75" swimtime="00:00:37.65" resultid="42123" heatid="45027" lane="7" entrytime="00:00:37.10" entrycourse="LCM" />
                <RESULT eventid="2430" points="693" reactiontime="+95" swimtime="00:00:31.38" resultid="42124" heatid="45071" lane="5" entrytime="00:00:32.49" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filipe Teixeira" lastname="Sa" birthdate="1978-10-31" gender="M" nation="POR" license="206936" swrid="5277962" athleteid="42187">
              <RESULTS>
                <RESULT comment="722 - Tocou com uma mão na parede na viragem aos 150 m - SW 7.6" eventid="2622" reactiontime="+104" status="DSQ" swimtime="00:03:15.20" resultid="42188" heatid="44878" lane="6" entrytime="00:03:10.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.31" />
                    <SPLIT distance="100" swimtime="00:01:29.28" />
                    <SPLIT distance="150" swimtime="00:02:21.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="456" reactiontime="+82" swimtime="00:00:33.63" resultid="42189" heatid="44896" lane="6" entrytime="00:00:36.16" entrycourse="LCM" />
                <RESULT eventid="2188" points="543" reactiontime="+84" swimtime="00:00:37.39" resultid="42190" heatid="44948" lane="5" entrytime="00:00:37.39" entrycourse="LCM" />
                <RESULT eventid="2385" points="365" reactiontime="+80" swimtime="00:03:05.20" resultid="42191" heatid="44975" lane="7" entrytime="00:06:33.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.97" />
                    <SPLIT distance="100" swimtime="00:01:30.04" />
                    <SPLIT distance="150" swimtime="00:02:22.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="507" reactiontime="+90" swimtime="00:01:26.08" resultid="42192" heatid="44998" lane="8" entrytime="00:01:25.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Fernanda" lastname="Goncalves" birthdate="1966-03-01" gender="F" nation="POR" license="117412" swrid="4496936" athleteid="42137">
              <RESULTS>
                <RESULT eventid="2203" status="DNS" swimtime="00:00:00.00" resultid="42138" heatid="44882" lane="6" entrytime="00:01:34.15" entrycourse="LCM" />
                <RESULT eventid="2278" points="524" reactiontime="+99" swimtime="00:02:53.31" resultid="42139" heatid="44904" lane="8" entrytime="00:03:07.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:01:21.59" />
                    <SPLIT distance="150" swimtime="00:02:07.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="600" reactiontime="+91" swimtime="00:01:15.47" resultid="42140" heatid="44956" lane="7" entrytime="00:01:16.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="605" reactiontime="+76" swimtime="00:00:42.26" resultid="42141" heatid="45026" lane="2" entrytime="00:00:41.29" entrycourse="LCM" />
                <RESULT eventid="2430" points="676" reactiontime="+95" swimtime="00:00:33.73" resultid="42142" heatid="45071" lane="8" entrytime="00:00:34.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Celso Fernando" lastname="Ribeiro" birthdate="1969-07-23" gender="M" nation="POR" license="127787" swrid="4905842" athleteid="42178">
              <RESULTS>
                <RESULT eventid="1058" points="405" swimtime="00:12:24.77" resultid="42179" heatid="45083" lane="5" entrytime="00:12:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.77" />
                    <SPLIT distance="200" swimtime="00:03:03.27" />
                    <SPLIT distance="300" swimtime="00:04:38.03" />
                    <SPLIT distance="400" swimtime="00:06:13.52" />
                    <SPLIT distance="500" swimtime="00:07:47.25" />
                    <SPLIT distance="600" swimtime="00:09:21.56" />
                    <SPLIT distance="700" swimtime="00:10:56.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="493" reactiontime="+75" swimtime="00:02:41.02" resultid="42180" heatid="45092" lane="1" entrytime="00:03:03.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:18.04" />
                    <SPLIT distance="150" swimtime="00:02:00.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="432" reactiontime="+72" swimtime="00:03:10.65" resultid="42181" heatid="44978" lane="3" entrytime="00:03:09.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                    <SPLIT distance="100" swimtime="00:01:31.89" />
                    <SPLIT distance="150" swimtime="00:02:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" points="351" reactiontime="+72" swimtime="00:03:28.44" resultid="42182" heatid="45029" lane="5" entrytime="00:03:16.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.64" />
                    <SPLIT distance="100" swimtime="00:01:42.35" />
                    <SPLIT distance="150" swimtime="00:02:35.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="431" reactiontime="+73" swimtime="00:06:59.92" resultid="42183" heatid="45060" lane="2" entrytime="00:06:42.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.42" />
                    <SPLIT distance="100" swimtime="00:01:38.18" />
                    <SPLIT distance="150" swimtime="00:02:34.73" />
                    <SPLIT distance="200" swimtime="00:03:32.03" />
                    <SPLIT distance="250" swimtime="00:04:34.54" />
                    <SPLIT distance="300" swimtime="00:05:34.96" />
                    <SPLIT distance="350" swimtime="00:06:21.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joana Aguiar" lastname="Rodrigues" birthdate="1993-02-03" gender="F" nation="POR" license="15401" swrid="4061190" athleteid="42184">
              <RESULTS>
                <RESULT eventid="2607" points="494" reactiontime="+81" swimtime="00:00:41.28" resultid="42185" heatid="45102" lane="4" entrytime="00:00:41.98" entrycourse="LCM" />
                <RESULT eventid="2430" points="690" reactiontime="+75" swimtime="00:00:29.53" resultid="42186" heatid="45073" lane="3" entrytime="00:00:29.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alfredo Gouveia" lastname="Ferraria" birthdate="1957-06-07" gender="M" nation="POR" license="102458" swrid="4840961" athleteid="42125">
              <RESULTS>
                <RESULT eventid="2622" points="114" swimtime="00:05:51.24" resultid="42126" heatid="44872" lane="5" entrytime="00:05:24.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.18" />
                    <SPLIT distance="100" swimtime="00:02:51.77" />
                    <SPLIT distance="150" swimtime="00:04:23.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="123" reactiontime="+105" swimtime="00:01:07.55" resultid="42127" heatid="44939" lane="8" entrytime="00:01:00.64" entrycourse="LCM" />
                <RESULT eventid="2293" points="79" reactiontime="+74" swimtime="00:01:16.66" resultid="42128" heatid="45014" lane="1" entrytime="00:01:11.29" entrycourse="LCM" />
                <RESULT eventid="2445" points="112" reactiontime="+132" swimtime="00:02:39.69" resultid="42129" heatid="44990" lane="3" entrytime="00:02:25.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="134" reactiontime="+116" swimtime="00:00:53.28" resultid="42130" heatid="45033" lane="3" entrytime="00:00:52.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cristian" lastname="Aita" birthdate="1977-11-03" gender="M" nation="POR" license="213924" swrid="5464030" athleteid="42063">
              <RESULTS>
                <RESULT eventid="1058" points="347" swimtime="00:12:28.59" resultid="42064" heatid="45084" lane="1" entrytime="00:12:03.36">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.97" />
                    <SPLIT distance="200" swimtime="00:02:51.99" />
                    <SPLIT distance="300" swimtime="00:04:24.57" />
                    <SPLIT distance="400" swimtime="00:06:00.57" />
                    <SPLIT distance="500" swimtime="00:07:38.51" />
                    <SPLIT distance="600" swimtime="00:09:16.56" />
                    <SPLIT distance="700" swimtime="00:10:53.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2622" points="411" reactiontime="+85" swimtime="00:03:22.81" resultid="42065" heatid="44876" lane="4" entrytime="00:03:25.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.84" />
                    <SPLIT distance="100" swimtime="00:01:37.52" />
                    <SPLIT distance="150" swimtime="00:02:31.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" status="DNS" swimtime="00:00:00.00" resultid="42066" heatid="44978" lane="5" entrytime="00:03:09.52" />
                <RESULT eventid="2263" points="343" reactiontime="+82" swimtime="00:06:03.22" resultid="42067" heatid="45130" lane="8" entrytime="00:05:35.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:01:18.09" />
                    <SPLIT distance="150" swimtime="00:02:01.12" />
                    <SPLIT distance="200" swimtime="00:02:45.89" />
                    <SPLIT distance="250" swimtime="00:03:33.56" />
                    <SPLIT distance="300" swimtime="00:04:21.93" />
                    <SPLIT distance="350" swimtime="00:05:12.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="411" reactiontime="+76" swimtime="00:00:38.17" resultid="42068" heatid="45019" lane="1" entrytime="00:00:39.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Fernando" lastname="Sousa" birthdate="1965-08-16" gender="M" nation="POR" license="202718" swrid="4845984" athleteid="42222">
              <RESULTS>
                <RESULT eventid="2622" points="621" reactiontime="+76" swimtime="00:03:11.55" resultid="42223" heatid="44878" lane="7" entrytime="00:03:14.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                    <SPLIT distance="100" swimtime="00:01:31.65" />
                    <SPLIT distance="150" swimtime="00:02:21.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2537" points="555" reactiontime="+67" swimtime="00:01:23.06" resultid="42224" heatid="44887" lane="6" entrytime="00:01:24.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="571" reactiontime="+78" swimtime="00:03:01.93" resultid="42225" heatid="44919" lane="4" entrytime="00:03:10.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.29" />
                    <SPLIT distance="100" swimtime="00:01:31.69" />
                    <SPLIT distance="150" swimtime="00:02:19.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="650" reactiontime="+107" swimtime="00:00:36.14" resultid="42226" heatid="45019" lane="5" entrytime="00:00:37.33" entrycourse="LCM" />
                <RESULT eventid="2445" points="598" reactiontime="+83" swimtime="00:01:26.22" resultid="42227" heatid="44997" lane="5" entrytime="00:01:26.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carla Santa" lastname="Barbara" birthdate="1975-03-22" gender="F" nation="POR" license="118948" swrid="4590248" athleteid="42081">
              <RESULTS>
                <RESULT comment="Rec Nac Esc E" eventid="2278" points="707" reactiontime="+81" swimtime="00:02:29.60" resultid="42082" heatid="44905" lane="6" entrytime="00:02:25.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                    <SPLIT distance="100" swimtime="00:01:11.90" />
                    <SPLIT distance="150" swimtime="00:01:51.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="645" reactiontime="+75" swimtime="00:00:41.89" resultid="42083" heatid="45103" lane="8" entrytime="00:00:41.73" entrycourse="LCM" />
                <RESULT eventid="2637" points="713" reactiontime="+75" swimtime="00:01:07.08" resultid="42084" heatid="44957" lane="3" entrytime="00:01:06.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="729" reactiontime="+75" swimtime="00:00:30.85" resultid="42085" heatid="45072" lane="4" entrytime="00:00:30.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alfredo Coelho" lastname="Magalhaes" birthdate="1953-11-29" gender="M" nation="POR" license="210499" swrid="5365300" athleteid="42149">
              <RESULTS>
                <RESULT eventid="2622" points="282" swimtime="00:04:45.76" resultid="42150" heatid="44873" lane="7" entrytime="00:04:54.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.38" />
                    <SPLIT distance="100" swimtime="00:02:20.44" />
                    <SPLIT distance="150" swimtime="00:03:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="94" reactiontime="+104" swimtime="00:05:53.01" resultid="42151" heatid="44917" lane="8" entrytime="00:04:35.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.68" />
                    <SPLIT distance="100" swimtime="00:02:51.89" />
                    <SPLIT distance="150" swimtime="00:04:26.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="188" swimtime="00:01:00.19" resultid="42152" heatid="44938" lane="3" entrytime="00:01:01.37" entrycourse="LCM" />
                <RESULT eventid="2293" points="126" reactiontime="+90" swimtime="00:01:06.81" resultid="42153" heatid="45014" lane="2" entrytime="00:01:09.26" entrycourse="LCM" />
                <RESULT eventid="2445" points="252" swimtime="00:02:10.38" resultid="42154" heatid="44991" lane="7" entrytime="00:02:15.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia Manso" lastname="Marchioro" birthdate="1993-03-08" gender="F" nation="ITA" license="213958" swrid="5464031" athleteid="42155">
              <RESULTS>
                <RESULT eventid="2203" points="478" reactiontime="+66" swimtime="00:01:25.03" resultid="42156" heatid="44882" lane="5" entrytime="00:01:32.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2308" points="433" reactiontime="+87" swimtime="00:03:13.05" resultid="42157" heatid="44915" lane="3" entrytime="00:02:25.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                    <SPLIT distance="100" swimtime="00:01:29.86" />
                    <SPLIT distance="150" swimtime="00:02:21.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="377" reactiontime="+82" swimtime="00:01:19.22" resultid="42158" heatid="44956" lane="5" entrytime="00:01:13.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="500" reactiontime="+92" swimtime="00:00:38.51" resultid="42159" heatid="45026" lane="5" entrytime="00:00:39.12" entrycourse="LCM" />
                <RESULT eventid="2430" points="431" reactiontime="+81" swimtime="00:00:34.55" resultid="42160" heatid="45070" lane="3" entrytime="00:00:35.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Pedro" lastname="Soares" birthdate="1967-08-29" gender="M" nation="POR" license="130450" swrid="4995541" athleteid="42216">
              <RESULTS>
                <RESULT eventid="2537" points="620" reactiontime="+99" swimtime="00:01:17.20" resultid="42217" heatid="44887" lane="3" entrytime="00:01:19.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="596" reactiontime="+64" swimtime="00:02:56.24" resultid="42218" heatid="44921" lane="5" entrytime="00:02:20.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.71" />
                    <SPLIT distance="100" swimtime="00:01:28.71" />
                    <SPLIT distance="150" swimtime="00:02:14.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="704" reactiontime="+84" swimtime="00:01:03.90" resultid="42219" heatid="45113" lane="3" entrytime="00:01:03.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="828" reactiontime="+62" swimtime="00:00:31.69" resultid="42220" heatid="45022" lane="6" entrytime="00:00:31.13" entrycourse="LCM" />
                <RESULT eventid="2652" points="755" reactiontime="+80" swimtime="00:00:27.58" resultid="42221" heatid="45045" lane="4" entrytime="00:00:27.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo Monteiro" lastname="Pinto" birthdate="1964-03-26" gender="M" nation="POR" license="211230" swrid="5425459" athleteid="42164">
              <RESULTS>
                <RESULT comment="603 - Após viragem saiu em posição ventral aos 150 m - SW 6.2" eventid="2218" reactiontime="+106" status="DSQ" swimtime="00:05:10.87" resultid="42165" heatid="44917" lane="1" entrytime="00:04:35.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.97" />
                    <SPLIT distance="100" swimtime="00:02:29.12" />
                    <SPLIT distance="150" swimtime="00:03:49.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="136" reactiontime="+139" swimtime="00:01:00.25" resultid="42166" heatid="44938" lane="2" entrytime="00:01:03.37" />
                <RESULT eventid="2263" points="159" reactiontime="+128" swimtime="00:08:29.30" resultid="42167" heatid="45124" lane="4" entrytime="00:08:17.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.89" />
                    <SPLIT distance="100" swimtime="00:01:53.31" />
                    <SPLIT distance="150" swimtime="00:02:58.41" />
                    <SPLIT distance="200" swimtime="00:04:04.62" />
                    <SPLIT distance="250" swimtime="00:05:11.08" />
                    <SPLIT distance="300" swimtime="00:06:19.29" />
                    <SPLIT distance="350" swimtime="00:07:27.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="101" reactiontime="+101" swimtime="00:01:07.20" resultid="42168" heatid="45014" lane="6" entrytime="00:01:07.83" entrycourse="LCM" />
                <RESULT eventid="2445" points="159" reactiontime="+122" swimtime="00:02:14.02" resultid="42169" heatid="44991" lane="8" entrytime="00:02:16.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Celso Ruben" lastname="Barbosa" birthdate="1977-10-09" gender="M" nation="POR" license="201888" swrid="5187807" athleteid="42086">
              <RESULTS>
                <RESULT eventid="2507" points="662" reactiontime="+71" swimtime="00:02:15.93" resultid="42087" heatid="45096" lane="2" entrytime="00:02:13.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                    <SPLIT distance="100" swimtime="00:01:08.10" />
                    <SPLIT distance="150" swimtime="00:01:42.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2323" points="564" reactiontime="+73" swimtime="00:01:11.02" resultid="42088" heatid="44929" lane="7" entrytime="00:01:08.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="588" reactiontime="+83" swimtime="00:05:03.51" resultid="42089" heatid="45131" lane="8" entrytime="00:05:17.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:01:12.83" />
                    <SPLIT distance="150" swimtime="00:01:52.12" />
                    <SPLIT distance="200" swimtime="00:02:32.16" />
                    <SPLIT distance="250" swimtime="00:03:11.87" />
                    <SPLIT distance="300" swimtime="00:03:50.57" />
                    <SPLIT distance="350" swimtime="00:04:27.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" points="324" reactiontime="+81" swimtime="00:03:12.59" resultid="42090" heatid="45030" lane="1" entrytime="00:03:05.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.03" />
                    <SPLIT distance="100" swimtime="00:01:35.48" />
                    <SPLIT distance="150" swimtime="00:02:27.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="698" reactiontime="+74" swimtime="00:00:27.70" resultid="42091" heatid="45046" lane="5" entrytime="00:00:27.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hugo Miguel" lastname="Vilas" birthdate="1978-11-02" gender="M" nation="POR" license="211227" swrid="4780256" athleteid="42245">
              <RESULTS>
                <RESULT eventid="2537" status="DNS" swimtime="00:00:00.00" resultid="42246" heatid="44888" lane="6" entrytime="00:01:13.36" />
                <RESULT eventid="2415" points="362" reactiontime="+83" swimtime="00:01:16.17" resultid="42247" heatid="45106" lane="6" entrytime="00:01:27.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="328" reactiontime="+66" swimtime="00:00:41.17" resultid="42248" heatid="45019" lane="6" entrytime="00:00:37.76" />
                <RESULT eventid="2652" points="454" reactiontime="+80" swimtime="00:00:31.96" resultid="42249" heatid="45041" lane="8" entrytime="00:00:31.53" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia Isabel" lastname="Pereira" birthdate="1981-01-19" gender="F" nation="POR" license="106652" swrid="4507633" athleteid="42161">
              <RESULTS>
                <RESULT eventid="2607" points="433" reactiontime="+83" swimtime="00:00:46.19" resultid="42162" heatid="45102" lane="8" entrytime="00:00:44.25" entrycourse="LCM" />
                <RESULT eventid="2430" points="467" reactiontime="+80" swimtime="00:00:35.36" resultid="42163" heatid="45069" lane="1" entrytime="00:00:38.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Nuno" lastname="Pires" birthdate="1975-03-04" gender="M" nation="POR" license="210671" swrid="5371327" athleteid="42170">
              <RESULTS>
                <RESULT eventid="2682" points="320" reactiontime="+88" swimtime="00:00:38.83" resultid="42171" heatid="44895" lane="8" entrytime="00:00:40.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Joao" lastname="Taborda" birthdate="1967-10-22" gender="F" nation="POR" license="123373" swrid="4756614" athleteid="42240">
              <RESULTS>
                <RESULT eventid="2173" points="406" swimtime="00:04:07.35" resultid="42241" heatid="45088" lane="6" entrytime="00:03:53.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.39" />
                    <SPLIT distance="100" swimtime="00:01:58.88" />
                    <SPLIT distance="150" swimtime="00:03:03.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="351" reactiontime="+100" swimtime="00:00:52.02" resultid="42242" heatid="45100" lane="6" entrytime="00:00:49.82" entrycourse="LCM" />
                <RESULT eventid="2460" points="378" reactiontime="+104" swimtime="00:01:54.82" resultid="42243" heatid="45120" lane="5" entrytime="00:01:50.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="255" reactiontime="+107" swimtime="00:00:44.77" resultid="42244" heatid="45067" lane="7" entrytime="00:00:46.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Marcos" lastname="Madureira" birthdate="1964-04-25" gender="M" nation="POR" license="207162" swrid="5282675" athleteid="42143">
              <RESULTS>
                <RESULT eventid="2622" points="324" reactiontime="+103" swimtime="00:03:57.82" resultid="42144" heatid="44876" lane="5" entrytime="00:03:25.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.99" />
                    <SPLIT distance="100" swimtime="00:01:57.02" />
                    <SPLIT distance="150" swimtime="00:03:01.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="330" reactiontime="+101" swimtime="00:00:44.90" resultid="42145" heatid="44944" lane="1" entrytime="00:00:44.29" entrycourse="LCM" />
                <RESULT eventid="2415" points="346" reactiontime="+94" swimtime="00:01:25.55" resultid="42146" heatid="45114" lane="8" entrytime="00:01:03.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="346" reactiontime="+93" swimtime="00:01:43.40" resultid="42147" heatid="44994" lane="3" entrytime="00:01:43.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="392" reactiontime="+97" swimtime="00:00:36.33" resultid="42148" heatid="45037" lane="2" entrytime="00:00:35.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carla Sofia" lastname="Santos" birthdate="1989-04-07" gender="F" nation="POR" license="204832" swrid="5215226" athleteid="42199">
              <RESULTS>
                <RESULT eventid="2338" status="DNS" swimtime="00:00:00.00" resultid="42200" heatid="44892" lane="6" entrytime="00:00:32.59" entrycourse="LCM" />
                <RESULT eventid="2278" status="DNS" swimtime="00:00:00.00" resultid="42201" heatid="44905" lane="7" entrytime="00:02:36.05" />
                <RESULT eventid="2637" points="531" reactiontime="+61" swimtime="00:01:11.93" resultid="42202" heatid="44957" lane="7" entrytime="00:01:09.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="587" reactiontime="+74" swimtime="00:00:31.59" resultid="42203" heatid="45072" lane="5" entrytime="00:00:30.47" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Catarina Matos" lastname="Araujo" birthdate="1991-05-31" gender="F" nation="POR" license="15403" swrid="4574374" athleteid="42075">
              <RESULTS>
                <RESULT eventid="2338" points="454" reactiontime="+95" swimtime="00:00:37.21" resultid="42076" heatid="44891" lane="5" entrytime="00:00:36.28" entrycourse="LCM" />
                <RESULT eventid="2278" points="335" reactiontime="+95" swimtime="00:03:03.46" resultid="42077" heatid="44904" lane="6" entrytime="00:03:02.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                    <SPLIT distance="100" swimtime="00:01:25.51" />
                    <SPLIT distance="150" swimtime="00:02:14.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2552" points="258" reactiontime="+90" swimtime="00:01:41.32" resultid="42078" heatid="44923" lane="7" entrytime="00:01:59.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="377" reactiontime="+98" swimtime="00:01:20.62" resultid="42079" heatid="44956" lane="2" entrytime="00:01:16.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="461" reactiontime="+91" swimtime="00:00:34.25" resultid="42080" heatid="45071" lane="2" entrytime="00:00:33.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vivien Patricia" lastname="Silva" birthdate="1962-12-08" gender="F" nation="BRA" license="212365" athleteid="42204">
              <RESULTS>
                <RESULT eventid="2203" points="336" reactiontime="+87" swimtime="00:01:52.37" resultid="42205" heatid="44881" lane="4" entrytime="00:01:45.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2338" points="321" reactiontime="+97" swimtime="00:00:46.44" resultid="42206" heatid="44890" lane="2" entrytime="00:00:46.99" entrycourse="LCM" />
                <RESULT eventid="2308" points="347" reactiontime="+83" swimtime="00:03:57.60" resultid="42207" heatid="44915" lane="2" entrytime="00:02:36.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.32" />
                    <SPLIT distance="100" swimtime="00:01:57.44" />
                    <SPLIT distance="150" swimtime="00:02:57.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="316" reactiontime="+96" swimtime="00:07:06.87" resultid="42208" heatid="45010" lane="6" entrytime="00:07:19.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.33" />
                    <SPLIT distance="100" swimtime="00:01:40.47" />
                    <SPLIT distance="150" swimtime="00:02:33.81" />
                    <SPLIT distance="200" swimtime="00:03:29.10" />
                    <SPLIT distance="250" swimtime="00:04:23.05" />
                    <SPLIT distance="300" swimtime="00:05:18.16" />
                    <SPLIT distance="350" swimtime="00:06:12.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="304" reactiontime="+86" swimtime="00:00:53.16" resultid="42209" heatid="45024" lane="6" entrytime="00:00:51.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Alexandre" lastname="Sousa" birthdate="1982-04-09" gender="M" nation="POR" license="123374" swrid="4756745" athleteid="42228">
              <RESULTS>
                <RESULT eventid="2622" points="643" reactiontime="+74" swimtime="00:02:55.32" resultid="42229" heatid="44879" lane="8" entrytime="00:02:54.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                    <SPLIT distance="100" swimtime="00:01:25.50" />
                    <SPLIT distance="150" swimtime="00:02:11.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="688" reactiontime="+71" swimtime="00:00:28.90" resultid="42230" heatid="44900" lane="8" entrytime="00:00:29.74" entrycourse="LCM" />
                <RESULT eventid="2323" status="DNS" swimtime="00:00:00.00" resultid="42231" heatid="44930" lane="5" entrytime="00:00:59.36" />
                <RESULT eventid="2188" points="586" reactiontime="+68" swimtime="00:00:34.90" resultid="42232" heatid="44949" lane="6" entrytime="00:00:35.29" entrycourse="LCM" />
                <RESULT eventid="2445" points="611" reactiontime="+69" swimtime="00:01:18.31" resultid="42233" heatid="44999" lane="8" entrytime="00:01:18.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno Miguel" lastname="Santos" birthdate="1976-07-27" gender="M" nation="POR" license="14631" swrid="4575729" athleteid="42193">
              <RESULTS>
                <RESULT eventid="2537" points="574" reactiontime="+99" swimtime="00:01:14.42" resultid="42194" heatid="44888" lane="1" entrytime="00:01:16.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="711" reactiontime="+70" swimtime="00:00:29.75" resultid="42195" heatid="44899" lane="3" entrytime="00:00:30.30" entrycourse="LCM" />
                <RESULT eventid="2507" points="580" reactiontime="+77" swimtime="00:02:23.13" resultid="42196" heatid="45095" lane="6" entrytime="00:02:22.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:10.26" />
                    <SPLIT distance="150" swimtime="00:01:47.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="456" reactiontime="+75" swimtime="00:02:56.20" resultid="42197" heatid="44920" lane="4" entrytime="00:02:50.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:23.26" />
                    <SPLIT distance="150" swimtime="00:02:09.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2323" points="626" reactiontime="+78" swimtime="00:01:10.62" resultid="42198" heatid="44928" lane="5" entrytime="00:01:09.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Tiago" lastname="Soares" birthdate="1970-07-18" gender="M" nation="POR" license="201938" swrid="5191965" athleteid="42210">
              <RESULTS>
                <RESULT eventid="2622" points="416" reactiontime="+86" swimtime="00:03:34.26" resultid="42211" heatid="44876" lane="3" entrytime="00:03:25.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.74" />
                    <SPLIT distance="100" swimtime="00:01:45.34" />
                    <SPLIT distance="150" swimtime="00:02:42.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="437" reactiontime="+88" swimtime="00:00:36.40" resultid="42212" heatid="44894" lane="5" entrytime="00:00:41.30" />
                <RESULT eventid="2188" points="466" reactiontime="+78" swimtime="00:00:40.13" resultid="42213" heatid="44947" lane="1" entrytime="00:00:39.34" entrycourse="LCM" />
                <RESULT eventid="2445" points="477" reactiontime="+77" swimtime="00:01:32.73" resultid="42214" heatid="44996" lane="2" entrytime="00:01:33.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="486" reactiontime="+80" swimtime="00:00:31.94" resultid="42215" heatid="45040" lane="6" entrytime="00:00:31.91" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Aderito" lastname="Chaves" birthdate="1970-10-30" gender="M" nation="POR" license="127786" swrid="4905840" athleteid="42108">
              <RESULTS>
                <RESULT eventid="2537" status="DNS" swimtime="00:00:00.00" resultid="42109" heatid="44888" lane="3" entrytime="00:01:11.70" entrycourse="LCM" />
                <RESULT eventid="2507" status="DNS" swimtime="00:00:00.00" resultid="42110" heatid="45096" lane="1" entrytime="00:02:16.15" />
                <RESULT eventid="2218" status="DNS" swimtime="00:00:00.00" resultid="42111" heatid="44921" lane="1" entrytime="00:02:42.23" entrycourse="LCM" />
                <RESULT eventid="2293" status="DNS" swimtime="00:00:00.00" resultid="42112" heatid="45022" lane="1" entrytime="00:00:32.63" entrycourse="LCM" />
                <RESULT eventid="2248" status="DNS" swimtime="00:00:00.00" resultid="42113" heatid="45062" lane="8" entrytime="00:05:45.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo Jorge" lastname="Cohen" birthdate="1959-08-22" gender="M" nation="POR" license="26838" swrid="4319462" athleteid="42114">
              <RESULTS>
                <RESULT eventid="2682" points="443" reactiontime="+100" swimtime="00:00:38.18" resultid="42115" heatid="44894" lane="3" entrytime="00:00:41.30" entrycourse="LCM" />
                <RESULT eventid="2415" points="494" reactiontime="+103" swimtime="00:01:17.18" resultid="42116" heatid="45109" lane="7" entrytime="00:01:16.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="458" reactiontime="+82" swimtime="00:00:42.68" resultid="42117" heatid="45017" lane="3" entrytime="00:00:45.05" entrycourse="LCM" />
                <RESULT eventid="2652" points="601" reactiontime="+89" swimtime="00:00:32.37" resultid="42118" heatid="45040" lane="2" entrytime="00:00:31.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Margarida Bleck" lastname="Reis" birthdate="1968-01-22" gender="F" nation="POR" license="210540" swrid="5367932" athleteid="42172">
              <RESULTS>
                <RESULT eventid="1060" points="281" swimtime="00:15:03.52" resultid="42173" heatid="45077" lane="1" entrytime="00:14:17.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.10" />
                    <SPLIT distance="200" swimtime="00:03:37.15" />
                    <SPLIT distance="300" swimtime="00:05:33.27" />
                    <SPLIT distance="400" swimtime="00:07:29.73" />
                    <SPLIT distance="500" swimtime="00:09:25.54" />
                    <SPLIT distance="600" swimtime="00:11:20.58" />
                    <SPLIT distance="700" swimtime="00:13:14.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2338" points="270" reactiontime="+95" swimtime="00:00:46.76" resultid="42174" heatid="44890" lane="6" entrytime="00:00:46.31" entrycourse="LCM" />
                <RESULT eventid="2233" points="328" reactiontime="+108" swimtime="00:03:48.75" resultid="42175" heatid="44972" lane="6" entrytime="00:03:25.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.65" />
                    <SPLIT distance="100" swimtime="00:01:49.81" />
                    <SPLIT distance="150" swimtime="00:02:56.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="298" reactiontime="+90" swimtime="00:07:11.52" resultid="42176" heatid="45010" lane="4" entrytime="00:07:06.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.64" />
                    <SPLIT distance="100" swimtime="00:01:39.72" />
                    <SPLIT distance="150" swimtime="00:02:35.62" />
                    <SPLIT distance="200" swimtime="00:03:32.10" />
                    <SPLIT distance="250" swimtime="00:04:27.77" />
                    <SPLIT distance="300" swimtime="00:05:23.61" />
                    <SPLIT distance="350" swimtime="00:06:19.72" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="615 - Não efectuou movimento continuo e imediato na viragem aos 150 - SW 6.4" eventid="2400" status="DSQ" swimtime="00:00:00.00" resultid="42177" heatid="45063" lane="4" entrytime="00:08:22.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Teresa" lastname="Andrade" birthdate="1963-02-26" gender="F" nation="POR" license="203942" swrid="4174636" athleteid="42069">
              <RESULTS>
                <RESULT comment="709 - Movimento alternado de braços durante o percurso - SW 7.2" eventid="2173" status="DSQ" swimtime="00:03:36.32" resultid="42070" heatid="45089" lane="7" entrytime="00:03:32.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.92" />
                    <SPLIT distance="100" swimtime="00:01:41.86" />
                    <SPLIT distance="150" swimtime="00:02:38.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="661" reactiontime="+70" swimtime="00:00:43.39" resultid="42071" heatid="45102" lane="3" entrytime="00:00:42.77" entrycourse="LCM" />
                <RESULT eventid="2522" points="541" reactiontime="+75" swimtime="00:00:43.86" resultid="42072" heatid="45025" lane="3" entrytime="00:00:44.33" entrycourse="LCM" />
                <RESULT comment="Rec Nac Esc G" eventid="2460" points="665" reactiontime="+67" swimtime="00:01:37.10" resultid="42073" heatid="45122" lane="7" entrytime="00:01:38.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="612" reactiontime="+66" swimtime="00:00:34.86" resultid="42074" heatid="45071" lane="1" entrytime="00:00:34.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco Santos" lastname="Barros" birthdate="1972-03-17" gender="M" nation="POR" license="108661" swrid="4345381" athleteid="42092">
              <RESULTS>
                <RESULT eventid="1058" points="378" swimtime="00:12:12.92" resultid="42093" heatid="45084" lane="8" entrytime="00:12:03.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.12" />
                    <SPLIT distance="200" swimtime="00:02:53.36" />
                    <SPLIT distance="300" swimtime="00:04:27.13" />
                    <SPLIT distance="400" swimtime="00:06:01.83" />
                    <SPLIT distance="500" swimtime="00:07:36.00" />
                    <SPLIT distance="600" swimtime="00:09:09.59" />
                    <SPLIT distance="700" swimtime="00:10:43.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="384" reactiontime="+84" swimtime="00:02:44.16" resultid="42094" heatid="45094" lane="8" entrytime="00:02:39.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:16.74" />
                    <SPLIT distance="150" swimtime="00:02:00.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="397" reactiontime="+91" swimtime="00:05:48.47" resultid="42095" heatid="45129" lane="6" entrytime="00:05:48.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:01:20.23" />
                    <SPLIT distance="150" swimtime="00:02:04.96" />
                    <SPLIT distance="200" swimtime="00:02:49.45" />
                    <SPLIT distance="250" swimtime="00:03:34.40" />
                    <SPLIT distance="300" swimtime="00:04:20.23" />
                    <SPLIT distance="350" swimtime="00:05:05.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" points="273" reactiontime="+103" swimtime="00:03:34.62" resultid="42096" heatid="45029" lane="6" entrytime="00:03:25.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.54" />
                    <SPLIT distance="100" swimtime="00:01:44.75" />
                    <SPLIT distance="150" swimtime="00:02:39.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="373" reactiontime="+100" swimtime="00:07:00.01" resultid="42097" heatid="45060" lane="6" entrytime="00:06:42.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                    <SPLIT distance="100" swimtime="00:01:37.08" />
                    <SPLIT distance="150" swimtime="00:02:36.40" />
                    <SPLIT distance="200" swimtime="00:03:37.12" />
                    <SPLIT distance="250" swimtime="00:04:36.38" />
                    <SPLIT distance="300" swimtime="00:05:35.05" />
                    <SPLIT distance="350" swimtime="00:06:17.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Silvia Manuel" lastname="Sousa" birthdate="1984-10-24" gender="F" nation="POR" license="125537" swrid="5207467" athleteid="42234">
              <RESULTS>
                <RESULT eventid="2203" points="268" reactiontime="+76" swimtime="00:01:48.03" resultid="42235" heatid="44882" lane="4" entrytime="00:01:32.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2308" points="272" reactiontime="+89" swimtime="00:03:49.74" resultid="42236" heatid="44915" lane="5" entrytime="00:02:25.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.66" />
                    <SPLIT distance="100" swimtime="00:01:50.64" />
                    <SPLIT distance="150" swimtime="00:02:51.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="265" reactiontime="+88" swimtime="00:01:32.52" resultid="42237" heatid="44956" lane="3" entrytime="00:01:13.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="265" reactiontime="+90" swimtime="00:07:17.15" resultid="42238" heatid="45011" lane="6" entrytime="00:06:49.36">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.79" />
                    <SPLIT distance="100" swimtime="00:01:39.20" />
                    <SPLIT distance="150" swimtime="00:02:34.88" />
                    <SPLIT distance="200" swimtime="00:03:32.17" />
                    <SPLIT distance="250" swimtime="00:04:29.27" />
                    <SPLIT distance="300" swimtime="00:05:26.84" />
                    <SPLIT distance="350" swimtime="00:06:24.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="289" reactiontime="+86" swimtime="00:00:40.57" resultid="42239" heatid="45070" lane="5" entrytime="00:00:35.36" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CNN" nation="POR" region="ANL" clubid="41847" swrid="76748" name="Clube Nacional de Natacao" shortname="Nacional de Natacao">
          <ATHLETES>
            <ATHLETE firstname="Nuno Tiago" lastname="Varino" birthdate="1977-05-08" gender="M" nation="POR" license="210321" swrid="5350317" athleteid="41923">
              <RESULTS>
                <RESULT eventid="2415" points="573" reactiontime="+76" swimtime="00:01:05.40" resultid="41924" heatid="45112" lane="2" entrytime="00:01:05.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="403 - Falsa partida - SW 4.4" eventid="2652" reactiontime="+64" status="DSQ" swimtime="00:00:28.56" resultid="41925" heatid="45044" lane="7" entrytime="00:00:28.75" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PDEM" nation="POR" region="ANL" clubid="41767" swrid="66445" name="Palmela Desporto EEM" shortname="Palmela">
          <ATHLETES>
            <ATHLETE firstname="Andreia Azevedo" lastname="Almeida" birthdate="1986-04-04" gender="F" nation="POR" license="206080" swrid="5261578" athleteid="41768">
              <RESULTS>
                <RESULT comment="403 - Falsa partida - SW 4.4" eventid="2338" reactiontime="+81" status="DSQ" swimtime="00:01:02.41" resultid="41769" heatid="44889" lane="6" entrytime="00:01:04.33" entrycourse="LCM" />
                <RESULT eventid="2607" points="116" reactiontime="+125" swimtime="00:01:06.84" resultid="41770" heatid="45097" lane="3" entrytime="00:01:07.83" entrycourse="LCM" />
                <RESULT comment="804 - Braçada subaquática após a partida - SW 8.2" eventid="2233" reactiontime="+115" status="DSQ" swimtime="00:04:46.15" resultid="41771" heatid="44971" lane="6" entrytime="00:05:02.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.99" />
                    <SPLIT distance="100" swimtime="00:02:24.31" />
                    <SPLIT distance="150" swimtime="00:03:43.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="132" reactiontime="+105" swimtime="00:02:22.50" resultid="41772" heatid="45118" lane="7" entrytime="00:02:40.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="155" reactiontime="+109" swimtime="00:08:42.89" resultid="41773" heatid="45008" lane="5" entrytime="00:08:44.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.32" />
                    <SPLIT distance="100" swimtime="00:02:01.56" />
                    <SPLIT distance="150" swimtime="00:03:11.08" />
                    <SPLIT distance="200" swimtime="00:04:18.12" />
                    <SPLIT distance="250" swimtime="00:05:27.34" />
                    <SPLIT distance="300" swimtime="00:06:33.71" />
                    <SPLIT distance="350" swimtime="00:07:41.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="O2ADCP" nation="POR" region="ANALG" clubid="41760" swrid="85654" name="O2-Assoc. Desp. e Cult. de Portimao" shortname="O2 Portimao">
          <ATHLETES>
            <ATHLETE firstname="Manuel Edgar" lastname="Soares" birthdate="1954-07-24" gender="M" nation="POR" license="129129" swrid="4954912" athleteid="41761">
              <RESULTS>
                <RESULT eventid="2507" points="316" reactiontime="+92" swimtime="00:03:35.03" resultid="41762" heatid="45091" lane="2" entrytime="00:03:29.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                    <SPLIT distance="100" swimtime="00:01:38.12" />
                    <SPLIT distance="150" swimtime="00:02:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="357" reactiontime="+101" swimtime="00:00:48.64" resultid="41763" heatid="44940" lane="3" entrytime="00:00:50.40" entrycourse="LCM" />
                <RESULT eventid="2415" points="381" reactiontime="+88" swimtime="00:01:26.59" resultid="41764" heatid="45105" lane="4" entrytime="00:01:29.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="313" reactiontime="+93" swimtime="00:07:42.53" resultid="41765" heatid="45125" lane="2" entrytime="00:07:55.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.43" />
                    <SPLIT distance="100" swimtime="00:01:48.18" />
                    <SPLIT distance="150" swimtime="00:02:48.11" />
                    <SPLIT distance="200" swimtime="00:03:49.90" />
                    <SPLIT distance="250" swimtime="00:04:48.83" />
                    <SPLIT distance="300" swimtime="00:05:49.63" />
                    <SPLIT distance="350" swimtime="00:06:48.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="446" reactiontime="+94" swimtime="00:00:37.12" resultid="41766" heatid="45036" lane="5" entrytime="00:00:37.13" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CPCD" nation="POR" region="ANL" clubid="43804" swrid="76733" name="Centro Popular Cultura e Desporto" shortname="CPCD-Povoa St Iria">
          <ATHLETES>
            <ATHLETE firstname="Ana Rita" lastname="Lopes" birthdate="1992-08-07" gender="F" nation="POR" license="129056" swrid="5449809" athleteid="44027">
              <RESULTS>
                <RESULT eventid="2338" points="416" reactiontime="+89" swimtime="00:00:37.23" resultid="44028" heatid="44891" lane="2" entrytime="00:00:37.57" entrycourse="SCM" />
                <RESULT eventid="2552" points="303" reactiontime="+91" swimtime="00:01:32.38" resultid="44029" heatid="44923" lane="4" entrytime="00:01:31.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="401" reactiontime="+90" swimtime="00:03:13.32" resultid="44030" heatid="44973" lane="3" entrytime="00:03:10.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.60" />
                    <SPLIT distance="100" swimtime="00:01:36.43" />
                    <SPLIT distance="150" swimtime="00:02:29.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2667" points="321" reactiontime="+92" swimtime="00:03:26.59" resultid="44031" heatid="45031" lane="3" entrytime="00:03:24.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.58" />
                    <SPLIT distance="100" swimtime="00:01:36.53" />
                    <SPLIT distance="150" swimtime="00:02:31.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Fernando" lastname="Inacio" birthdate="1968-09-26" gender="M" nation="POR" license="213449" swrid="5449808" athleteid="44023">
              <RESULTS>
                <RESULT eventid="2682" points="324" reactiontime="+91" swimtime="00:00:40.23" resultid="44024" heatid="44895" lane="7" entrytime="00:00:40.05" entrycourse="SCM" />
                <RESULT eventid="2415" points="337" reactiontime="+101" swimtime="00:01:21.69" resultid="44025" heatid="45107" lane="6" entrytime="00:01:22.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="387" reactiontime="+105" swimtime="00:00:34.45" resultid="44026" heatid="45037" lane="3" entrytime="00:00:35.20" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nelson Duarte" lastname="Batista" birthdate="1980-01-31" gender="M" nation="POR" license="213084" swrid="4564487" athleteid="44017">
              <RESULTS>
                <RESULT eventid="2622" points="549" reactiontime="+99" swimtime="00:03:04.13" resultid="44018" heatid="44878" lane="5" entrytime="00:03:02.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                    <SPLIT distance="100" swimtime="00:01:26.80" />
                    <SPLIT distance="150" swimtime="00:02:15.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="467" reactiontime="+92" swimtime="00:00:33.37" resultid="44019" heatid="44897" lane="1" entrytime="00:00:34.96" />
                <RESULT eventid="2188" points="552" reactiontime="+85" swimtime="00:00:37.19" resultid="44020" heatid="44949" lane="8" entrytime="00:00:36.62" entrycourse="SCM" />
                <RESULT eventid="2445" points="554" reactiontime="+92" swimtime="00:01:23.57" resultid="44021" heatid="44998" lane="3" entrytime="00:01:20.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="444" reactiontime="+89" swimtime="00:00:32.20" resultid="44022" heatid="45041" lane="3" entrytime="00:00:30.94" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raquel Alexandra" lastname="Santos" birthdate="1995-11-15" gender="F" nation="POR" license="131722" athleteid="44032">
              <RESULTS>
                <RESULT eventid="2338" points="331" reactiontime="+86" swimtime="00:00:40.15" resultid="44033" heatid="44891" lane="6" entrytime="00:00:37.29" />
                <RESULT eventid="2552" points="257" reactiontime="+93" swimtime="00:01:37.63" resultid="44034" heatid="44924" lane="8" entrytime="00:01:30.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="408" reactiontime="+83" swimtime="00:03:12.10" resultid="44035" heatid="44973" lane="6" entrytime="00:03:11.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                    <SPLIT distance="100" swimtime="00:01:30.71" />
                    <SPLIT distance="150" swimtime="00:02:27.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2400" points="351" reactiontime="+87" swimtime="00:07:05.02" resultid="44036" heatid="45064" lane="2" entrytime="00:06:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.12" />
                    <SPLIT distance="100" swimtime="00:01:42.00" />
                    <SPLIT distance="150" swimtime="00:02:35.38" />
                    <SPLIT distance="200" swimtime="00:03:28.17" />
                    <SPLIT distance="250" swimtime="00:04:25.55" />
                    <SPLIT distance="300" swimtime="00:05:25.99" />
                    <SPLIT distance="350" swimtime="00:06:15.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="AAC" nation="POR" region="ANC" clubid="41848" swrid="68068" name="Associacao Academica de Coimbra" shortname="Academica de Coimbra">
          <ATHLETES>
            <ATHLETE firstname="Jose Manuel" lastname="Tojo" birthdate="1977-04-18" gender="M" nation="POR" license="112391" swrid="5220426" athleteid="41907">
              <RESULTS>
                <RESULT eventid="2537" points="375" reactiontime="+64" swimtime="00:01:25.08" resultid="41908" heatid="44886" lane="6" entrytime="00:01:34.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="389" reactiontime="+67" swimtime="00:03:03.37" resultid="41909" heatid="44919" lane="2" entrytime="00:03:17.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.34" />
                    <SPLIT distance="100" swimtime="00:01:29.60" />
                    <SPLIT distance="150" swimtime="00:02:17.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="437" reactiontime="+87" swimtime="00:02:54.44" resultid="41910" heatid="44979" lane="2" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                    <SPLIT distance="100" swimtime="00:01:25.31" />
                    <SPLIT distance="150" swimtime="00:02:15.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" points="276" reactiontime="+91" swimtime="00:03:23.16" resultid="41911" heatid="45029" lane="2" entrytime="00:03:31.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.69" />
                    <SPLIT distance="100" swimtime="00:01:33.08" />
                    <SPLIT distance="150" swimtime="00:02:27.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="388" reactiontime="+87" swimtime="00:06:27.88" resultid="41912" heatid="45060" lane="7" entrytime="00:06:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.83" />
                    <SPLIT distance="100" swimtime="00:01:28.75" />
                    <SPLIT distance="150" swimtime="00:02:23.06" />
                    <SPLIT distance="200" swimtime="00:03:15.61" />
                    <SPLIT distance="250" swimtime="00:04:11.86" />
                    <SPLIT distance="300" swimtime="00:05:07.37" />
                    <SPLIT distance="350" swimtime="00:05:49.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Isabel" lastname="Torres" birthdate="1960-03-26" gender="F" nation="POR" license="12229" swrid="4379334" athleteid="41913">
              <RESULTS>
                <RESULT eventid="2607" points="578" reactiontime="+106" swimtime="00:00:45.36" resultid="41914" heatid="45101" lane="3" entrytime="00:00:44.98" entrycourse="LCM" />
                <RESULT eventid="2637" points="520" reactiontime="+95" swimtime="00:01:27.40" resultid="41915" heatid="44954" lane="2" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="502" reactiontime="+94" swimtime="00:01:47.95" resultid="41916" heatid="45121" lane="6" entrytime="00:01:45.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="624" reactiontime="+92" swimtime="00:00:36.42" resultid="41917" heatid="45069" lane="4" entrytime="00:00:36.74" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nuno Avila" lastname="Franca" birthdate="1972-01-04" gender="M" nation="POR" license="153496" swrid="5119866" athleteid="41863">
              <RESULTS>
                <RESULT eventid="2622" points="364" reactiontime="+89" swimtime="00:03:35.27" resultid="41864" heatid="44876" lane="8" entrytime="00:03:35.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                    <SPLIT distance="100" swimtime="00:01:38.67" />
                    <SPLIT distance="150" swimtime="00:02:36.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2537" points="265" reactiontime="+78" swimtime="00:01:36.29" resultid="41865" heatid="44886" lane="4" entrytime="00:01:32.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="223" reactiontime="+78" swimtime="00:03:43.45" resultid="41866" heatid="44919" lane="1" entrytime="00:03:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.18" />
                    <SPLIT distance="100" swimtime="00:01:54.33" />
                    <SPLIT distance="150" swimtime="00:02:51.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="363" reactiontime="+83" swimtime="00:00:41.91" resultid="41867" heatid="44946" lane="7" entrytime="00:00:41.12" entrycourse="LCM" />
                <RESULT eventid="2445" points="368" reactiontime="+87" swimtime="00:01:36.15" resultid="41868" heatid="44995" lane="4" entrytime="00:01:35.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Virgilio Zacarias" lastname="Costa" birthdate="1931-07-21" gender="M" nation="POR" license="210706" swrid="5376435" athleteid="41849">
              <RESULTS>
                <RESULT eventid="2622" status="DNS" swimtime="00:00:00.00" resultid="41850" heatid="44872" lane="6" entrytime="00:06:18.23" entrycourse="LCM" />
                <RESULT eventid="2537" status="DNS" swimtime="00:00:00.00" resultid="41851" heatid="44884" lane="2" entrytime="00:04:00.00" />
                <RESULT eventid="2263" status="DNS" swimtime="00:00:00.00" resultid="41852" heatid="45124" lane="6" entrytime="00:10:00.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim Fidalgo" lastname="Freitas" birthdate="1947-04-16" gender="M" nation="POR" license="11231" swrid="4574902" athleteid="41869">
              <RESULTS>
                <RESULT eventid="2622" points="333" reactiontime="+137" swimtime="00:04:37.88" resultid="41870" heatid="44874" lane="5" entrytime="00:03:51.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.28" />
                    <SPLIT distance="100" swimtime="00:02:08.49" />
                    <SPLIT distance="150" swimtime="00:03:22.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="529" reactiontime="+123" swimtime="00:00:45.57" resultid="41871" heatid="44943" lane="4" entrytime="00:00:44.47" entrycourse="LCM" />
                <RESULT eventid="2445" points="443" reactiontime="+120" swimtime="00:01:52.34" resultid="41872" heatid="44993" lane="2" entrytime="00:01:48.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="276" reactiontime="+133" swimtime="00:00:53.58" resultid="41873" heatid="45015" lane="5" entrytime="00:00:55.90" entrycourse="LCM" />
                <RESULT eventid="2652" points="257" reactiontime="+121" swimtime="00:00:44.74" resultid="41874" heatid="45034" lane="6" entrytime="00:00:43.33" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marco Alexandre" lastname="Matos" birthdate="1982-11-18" gender="M" nation="POR" license="203815" swrid="4241889" athleteid="41875">
              <RESULTS>
                <RESULT eventid="2323" points="503" reactiontime="+82" swimtime="00:01:13.21" resultid="41876" heatid="44927" lane="8" entrytime="00:01:23.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="488" reactiontime="+77" swimtime="00:02:47.79" resultid="41877" heatid="44981" lane="8" entrytime="00:02:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:19.73" />
                    <SPLIT distance="150" swimtime="00:02:07.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="421" reactiontime="+76" swimtime="00:01:28.67" resultid="41878" heatid="44995" lane="2" entrytime="00:01:38.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="556" reactiontime="+81" swimtime="00:00:28.60" resultid="41879" heatid="45042" lane="7" entrytime="00:00:30.27" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco Jorge" lastname="Ferreira" birthdate="1962-04-08" gender="M" nation="POR" license="100124" swrid="4353016" athleteid="41857">
              <RESULTS>
                <RESULT eventid="2537" points="301" reactiontime="+75" swimtime="00:01:41.87" resultid="41858" heatid="44885" lane="4" entrytime="00:01:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="309" reactiontime="+84" swimtime="00:03:43.10" resultid="41859" heatid="44918" lane="4" entrytime="00:03:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.12" />
                    <SPLIT distance="100" swimtime="00:01:50.21" />
                    <SPLIT distance="150" swimtime="00:02:49.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="299" reactiontime="+109" swimtime="00:03:48.83" resultid="41860" heatid="44976" lane="5" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.53" />
                    <SPLIT distance="100" swimtime="00:01:50.51" />
                    <SPLIT distance="150" swimtime="00:03:02.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="277" reactiontime="+106" swimtime="00:07:03.66" resultid="41861" heatid="45127" lane="2" entrytime="00:06:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.89" />
                    <SPLIT distance="100" swimtime="00:01:40.33" />
                    <SPLIT distance="150" swimtime="00:02:35.12" />
                    <SPLIT distance="200" swimtime="00:03:29.93" />
                    <SPLIT distance="250" swimtime="00:04:24.52" />
                    <SPLIT distance="300" swimtime="00:05:19.09" />
                    <SPLIT distance="350" swimtime="00:06:12.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="340" reactiontime="+107" swimtime="00:00:38.11" resultid="41862" heatid="45037" lane="5" entrytime="00:00:35.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuel Monteiro" lastname="Tenreiro" birthdate="1940-06-03" gender="M" nation="POR" license="11175" swrid="4575953" athleteid="41903">
              <RESULTS>
                <RESULT eventid="2622" points="243" swimtime="00:05:51.88" resultid="41904" heatid="44872" lane="4" entrytime="00:05:22.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.71" />
                    <SPLIT distance="100" swimtime="00:02:59.65" />
                    <SPLIT distance="150" swimtime="00:04:30.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="301" reactiontime="+122" swimtime="00:01:05.34" resultid="41905" heatid="44938" lane="7" entrytime="00:01:07.67" entrycourse="LCM" />
                <RESULT eventid="2445" points="216" reactiontime="+147" swimtime="00:02:45.10" resultid="41906" heatid="44990" lane="7" entrytime="00:02:32.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:25.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eugenia Maria" lastname="Cunha" birthdate="1962-05-19" gender="F" nation="POR" license="26546" swrid="4574695" athleteid="41853">
              <RESULTS>
                <RESULT eventid="2338" points="496" reactiontime="+96" swimtime="00:00:40.21" resultid="41854" heatid="44891" lane="8" entrytime="00:00:39.15" entrycourse="LCM" />
                <RESULT eventid="2430" points="507" reactiontime="+77" swimtime="00:00:37.13" resultid="41855" heatid="45069" lane="7" entrytime="00:00:38.66" entrycourse="LCM" />
                <RESULT eventid="2552" status="DNS" swimtime="00:00:00.00" resultid="41856" heatid="44923" lane="5" entrytime="00:01:35.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabel Costa" lastname="Monteiro" birthdate="1953-01-28" gender="F" nation="POR" license="11174" swrid="4575287" athleteid="41880">
              <RESULTS>
                <RESULT eventid="2203" points="305" reactiontime="+103" swimtime="00:02:13.96" resultid="41881" heatid="44880" lane="7" entrytime="00:02:16.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="284" reactiontime="+102" swimtime="00:01:49.45" resultid="41882" heatid="44952" lane="4" entrytime="00:01:51.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="344" swimtime="00:00:57.96" resultid="41883" heatid="45023" lane="6" entrytime="00:01:04.93" entrycourse="LCM" />
                <RESULT eventid="2430" points="353" reactiontime="+114" swimtime="00:00:46.01" resultid="41884" heatid="45066" lane="3" entrytime="00:00:52.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Miguel" lastname="Tejo" birthdate="1969-05-30" gender="M" nation="POR" license="104306" swrid="4575950" athleteid="41897">
              <RESULTS>
                <RESULT eventid="2218" points="486" reactiontime="+95" swimtime="00:03:08.60" resultid="41898" heatid="44919" lane="5" entrytime="00:03:13.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.37" />
                    <SPLIT distance="100" swimtime="00:01:31.23" />
                    <SPLIT distance="150" swimtime="00:02:20.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="568" reactiontime="+99" swimtime="00:00:37.57" resultid="41899" heatid="44947" lane="6" entrytime="00:00:38.95" entrycourse="LCM" />
                <RESULT eventid="2385" points="489" reactiontime="+108" swimtime="00:03:03.02" resultid="41900" heatid="44979" lane="1" entrytime="00:03:00.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                    <SPLIT distance="100" swimtime="00:01:29.54" />
                    <SPLIT distance="150" swimtime="00:02:20.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="555" reactiontime="+101" swimtime="00:01:28.19" resultid="41901" heatid="44997" lane="1" entrytime="00:01:28.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="407" reactiontime="+101" swimtime="00:06:00.35" resultid="41902" heatid="45128" lane="4" entrytime="00:05:54.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:01:22.10" />
                    <SPLIT distance="150" swimtime="00:02:07.21" />
                    <SPLIT distance="200" swimtime="00:02:54.02" />
                    <SPLIT distance="250" swimtime="00:03:41.58" />
                    <SPLIT distance="300" swimtime="00:04:28.47" />
                    <SPLIT distance="350" swimtime="00:05:15.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Margarida" lastname="Urbano" birthdate="1963-03-01" gender="F" nation="POR" license="11355" swrid="4575970" athleteid="41918">
              <RESULTS>
                <RESULT eventid="2278" points="371" reactiontime="+103" swimtime="00:03:14.36" resultid="41919" heatid="44903" lane="3" entrytime="00:03:10.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.70" />
                    <SPLIT distance="100" swimtime="00:01:32.39" />
                    <SPLIT distance="150" swimtime="00:02:23.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="397" reactiontime="+98" swimtime="00:01:26.58" resultid="41920" heatid="44955" lane="7" entrytime="00:01:26.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="379" reactiontime="+96" swimtime="00:03:39.73" resultid="41921" heatid="44972" lane="7" entrytime="00:03:37.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.00" />
                    <SPLIT distance="100" swimtime="00:01:52.34" />
                    <SPLIT distance="150" swimtime="00:02:51.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="334" reactiontime="+115" swimtime="00:06:59.08" resultid="41922" heatid="45011" lane="2" entrytime="00:06:50.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.25" />
                    <SPLIT distance="100" swimtime="00:01:38.58" />
                    <SPLIT distance="150" swimtime="00:02:31.05" />
                    <SPLIT distance="200" swimtime="00:03:24.73" />
                    <SPLIT distance="250" swimtime="00:04:18.69" />
                    <SPLIT distance="300" swimtime="00:05:13.50" />
                    <SPLIT distance="350" swimtime="00:06:07.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Teresa" lastname="Oliveira" birthdate="1957-07-17" gender="F" nation="POR" license="10538" swrid="4575411" athleteid="41885">
              <RESULTS>
                <RESULT eventid="2203" points="201" reactiontime="+79" swimtime="00:02:21.16" resultid="41886" heatid="44880" lane="6" entrytime="00:02:10.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="383" reactiontime="+113" swimtime="00:00:52.01" resultid="41887" heatid="45099" lane="4" entrytime="00:00:50.97" entrycourse="LCM" />
                <RESULT eventid="2460" points="384" reactiontime="+122" swimtime="00:01:58.01" resultid="41888" heatid="45120" lane="7" entrytime="00:01:54.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="223" reactiontime="+86" swimtime="00:01:04.16" resultid="41889" heatid="45024" lane="8" entrytime="00:00:57.06" entrycourse="LCM" />
                <RESULT eventid="2430" points="287" reactiontime="+116" swimtime="00:00:47.19" resultid="41890" heatid="45068" lane="2" entrytime="00:00:42.26" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Manuel" lastname="Silva" birthdate="1964-01-20" gender="M" nation="POR" license="109826" swrid="4355906" athleteid="41891">
              <RESULTS>
                <RESULT eventid="2622" points="340" reactiontime="+108" swimtime="00:03:54.09" resultid="41892" heatid="44874" lane="4" entrytime="00:03:50.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.41" />
                    <SPLIT distance="100" swimtime="00:01:46.79" />
                    <SPLIT distance="150" swimtime="00:02:49.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2537" points="325" reactiontime="+94" swimtime="00:01:39.29" resultid="41893" heatid="44885" lane="3" entrytime="00:01:45.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="350" reactiontime="+101" swimtime="00:00:44.02" resultid="41894" heatid="44944" lane="7" entrytime="00:00:44.25" entrycourse="LCM" />
                <RESULT eventid="2445" points="355" reactiontime="+107" swimtime="00:01:42.53" resultid="41895" heatid="44993" lane="3" entrytime="00:01:45.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="337" reactiontime="+92" swimtime="00:00:44.95" resultid="41896" heatid="45017" lane="4" entrytime="00:00:44.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCCAM" nation="POR" region="ANMIN" clubid="42769" swrid="84575" name="Sporting Clube Caminhense" shortname="Sporting Caminhense">
          <ATHLETES>
            <ATHLETE firstname="Francisco Miguel" lastname="Vitoriano" birthdate="1971-05-23" gender="M" nation="POR" license="14397" swrid="4576019" athleteid="42790">
              <RESULTS>
                <RESULT eventid="2188" status="DNS" swimtime="00:00:00.00" resultid="42791" heatid="44947" lane="3" entrytime="00:00:38.65" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="42792" heatid="45041" lane="5" entrytime="00:00:30.84" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emilio Monteiro" lastname="Garmendia" birthdate="1982-09-30" gender="M" nation="POR" license="210558" swrid="5369506" athleteid="42770">
              <RESULTS>
                <RESULT eventid="2682" points="748" reactiontime="+74" swimtime="00:00:28.11" resultid="42771" heatid="44900" lane="5" entrytime="00:00:28.64" />
                <RESULT eventid="2415" points="719" reactiontime="+75" swimtime="00:00:58.01" resultid="42772" heatid="45116" lane="2" entrytime="00:00:57.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="776" reactiontime="+72" swimtime="00:00:25.60" resultid="42773" heatid="45048" lane="2" entrytime="00:00:25.92" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filipa Mendes" lastname="Pinheiro" birthdate="1992-06-27" gender="F" nation="POR" license="11056" swrid="4161354" athleteid="42781">
              <RESULTS>
                <RESULT eventid="2203" points="813" reactiontime="+62" swimtime="00:01:11.23" resultid="42782" heatid="44883" lane="4" entrytime="00:01:10.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2338" points="722" reactiontime="+73" swimtime="00:00:30.98" resultid="42783" heatid="44892" lane="5" entrytime="00:00:31.68" />
                <RESULT eventid="2308" points="758" reactiontime="+64" swimtime="00:02:40.22" resultid="42784" heatid="44915" lane="6" entrytime="00:02:36.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:01:16.61" />
                    <SPLIT distance="150" swimtime="00:01:58.43" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rec Nac Esc A" eventid="2522" points="873" reactiontime="+87" swimtime="00:00:31.98" resultid="42785" heatid="45027" lane="5" entrytime="00:00:33.27" />
                <RESULT eventid="2430" points="657" reactiontime="+70" swimtime="00:00:30.01" resultid="42786" heatid="45073" lane="7" entrytime="00:00:30.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique Mira" lastname="Godinho" birthdate="1988-07-29" gender="M" nation="POR" license="11664" swrid="4062840" athleteid="42777">
              <RESULTS>
                <RESULT eventid="2323" status="DNS" swimtime="00:00:00.00" resultid="42778" heatid="44929" lane="1" entrytime="00:01:08.73" />
                <RESULT eventid="2385" points="589" reactiontime="+84" swimtime="00:02:36.98" resultid="42779" heatid="44982" lane="1" entrytime="00:02:35.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:01:12.43" />
                    <SPLIT distance="150" swimtime="00:01:57.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="589" reactiontime="+89" swimtime="00:01:16.20" resultid="42780" heatid="44999" lane="2" entrytime="00:01:16.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andrea Helena" lastname="Pereira" birthdate="1977-02-13" gender="F" nation="POR" license="200630" swrid="4575470" athleteid="42774">
              <RESULTS>
                <RESULT eventid="2607" status="DNS" swimtime="00:00:00.00" resultid="42775" heatid="45098" lane="5" entrytime="00:00:56.93" />
                <RESULT eventid="2637" status="DNS" swimtime="00:00:00.00" resultid="42776" heatid="44953" lane="7" entrytime="00:01:46.29" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Alberto" lastname="Freixo" birthdate="1992-02-22" gender="M" nation="POR" license="11023" swrid="4269321" athleteid="42787">
              <RESULTS>
                <RESULT eventid="2218" status="DNS" swimtime="00:00:00.00" resultid="42788" heatid="44917" lane="4" entrytime="00:02:55.00" />
                <RESULT eventid="2293" status="DNS" swimtime="00:00:00.00" resultid="42789" heatid="45021" lane="3" entrytime="00:00:33.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SFGP" nation="POR" region="ANDS" clubid="41976" swrid="66448" name="Sociedade Filarmonica Gualdim Pais" shortname="Gualdim Pais">
          <ATHLETES>
            <ATHLETE firstname="Pedro Miguel" lastname="Caseiro" birthdate="1987-08-13" gender="M" nation="POR" license="212454" swrid="5424155" athleteid="41977">
              <RESULTS>
                <RESULT eventid="2323" points="320" reactiontime="+103" swimtime="00:01:22.87" resultid="41978" heatid="44927" lane="5" entrytime="00:01:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="410" reactiontime="+97" swimtime="00:01:08.41" resultid="41979" heatid="45110" lane="2" entrytime="00:01:11.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Miguel" lastname="Mesquita" birthdate="1989-05-23" gender="M" nation="POR" license="213362" swrid="4559308" athleteid="41984">
              <RESULTS>
                <RESULT eventid="2188" points="404" reactiontime="+89" swimtime="00:00:38.94" resultid="41985" heatid="44946" lane="3" entrytime="00:00:40.00" />
                <RESULT eventid="2415" points="428" reactiontime="+92" swimtime="00:01:07.42" resultid="41986" heatid="45112" lane="4" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo Jorge" lastname="Marques" birthdate="1986-08-22" gender="M" nation="POR" license="11495" swrid="4061332" athleteid="41980">
              <RESULTS>
                <RESULT eventid="2188" points="425" reactiontime="+86" swimtime="00:00:38.84" resultid="41981" heatid="44947" lane="5" entrytime="00:00:38.62" entrycourse="LCM" />
                <RESULT eventid="2415" points="526" reactiontime="+83" swimtime="00:01:04.39" resultid="41982" heatid="45114" lane="3" entrytime="00:01:01.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="429" reactiontime="+87" swimtime="00:02:55.06" resultid="41983" heatid="44980" lane="5" entrytime="00:02:49.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                    <SPLIT distance="100" swimtime="00:01:22.88" />
                    <SPLIT distance="150" swimtime="00:02:15.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CDF" nation="POR" region="ANCNP" clubid="42793" swrid="68061" name="Clube Desportivo Feirense" shortname="Feirense">
          <ATHLETES>
            <ATHLETE firstname="Hugo Gomes" lastname="Silva" birthdate="1994-09-10" gender="M" nation="POR" license="121434" swrid="4703325" athleteid="42864">
              <RESULTS>
                <RESULT eventid="2682" points="557" reactiontime="+67" swimtime="00:00:30.46" resultid="42865" heatid="44900" lane="6" entrytime="00:00:29.14" />
                <RESULT eventid="2323" points="465" reactiontime="+73" swimtime="00:01:13.37" resultid="42866" heatid="44928" lane="2" entrytime="00:01:11.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="420" reactiontime="+71" swimtime="00:01:09.02" resultid="42867" heatid="45113" lane="4" entrytime="00:01:03.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="428" reactiontime="+70" swimtime="00:02:47.16" resultid="42868" heatid="44980" lane="2" entrytime="00:02:53.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                    <SPLIT distance="100" swimtime="00:01:16.39" />
                    <SPLIT distance="150" swimtime="00:02:05.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="402" reactiontime="+70" swimtime="00:00:31.36" resultid="42869" heatid="45042" lane="3" entrytime="00:00:29.78" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabel Maria" lastname="Guimaraes" birthdate="1966-07-06" gender="F" nation="POR" license="204632" swrid="5207381" athleteid="42843">
              <RESULTS>
                <RESULT eventid="2607" points="210" reactiontime="+122" swimtime="00:01:03.51" resultid="42844" heatid="45097" lane="4" entrytime="00:01:05.05" entrycourse="LCM" />
                <RESULT eventid="2637" points="93" reactiontime="+102" swimtime="00:02:20.30" resultid="42845" heatid="44952" lane="8" entrytime="00:02:11.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mario Xavier" lastname="Rocha" birthdate="1970-12-13" gender="M" nation="POR" license="202205" swrid="4135956" athleteid="42860">
              <RESULTS>
                <RESULT eventid="2622" points="381" reactiontime="+102" swimtime="00:03:40.70" resultid="42861" heatid="44875" lane="3" entrytime="00:03:41.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.40" />
                    <SPLIT distance="100" swimtime="00:01:46.36" />
                    <SPLIT distance="150" swimtime="00:02:44.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="302" reactiontime="+93" swimtime="00:00:46.37" resultid="42862" heatid="44942" lane="7" entrytime="00:00:46.43" entrycourse="LCM" />
                <RESULT eventid="2445" points="366" reactiontime="+94" swimtime="00:01:41.26" resultid="42863" heatid="44994" lane="2" entrytime="00:01:43.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Gomes" lastname="Antoninho" birthdate="1978-10-20" gender="M" nation="POR" license="213338" swrid="5448808" athleteid="42800">
              <RESULTS>
                <RESULT eventid="2188" points="234" reactiontime="+87" swimtime="00:00:49.50" resultid="42801" heatid="44941" lane="5" entrytime="00:00:47.46" entrycourse="LCM" />
                <RESULT eventid="2415" points="199" reactiontime="+79" swimtime="00:01:32.94" resultid="42802" heatid="45106" lane="4" entrytime="00:01:26.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="245" reactiontime="+71" swimtime="00:01:49.63" resultid="42803" heatid="44993" lane="5" entrytime="00:01:45.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="222" reactiontime="+86" swimtime="00:00:46.88" resultid="42804" heatid="45016" lane="3" entrytime="00:00:50.04" />
                <RESULT eventid="2652" points="302" reactiontime="+81" swimtime="00:00:36.60" resultid="42805" heatid="45036" lane="4" entrytime="00:00:36.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Decio Manuel" lastname="Faria" birthdate="1972-06-30" gender="M" nation="POR" license="211173" swrid="5418290" athleteid="42827">
              <RESULTS>
                <RESULT eventid="2622" points="343" reactiontime="+95" swimtime="00:03:39.50" resultid="42828" heatid="44875" lane="2" entrytime="00:03:42.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.30" />
                    <SPLIT distance="100" swimtime="00:01:45.40" />
                    <SPLIT distance="150" swimtime="00:02:44.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="272" reactiontime="+99" swimtime="00:03:04.08" resultid="42829" heatid="45092" lane="3" entrytime="00:02:54.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                    <SPLIT distance="100" swimtime="00:01:25.09" />
                    <SPLIT distance="150" swimtime="00:02:15.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="248" reactiontime="+104" swimtime="00:00:45.79" resultid="42830" heatid="45016" lane="5" entrytime="00:00:48.97" />
                <RESULT eventid="2652" points="378" reactiontime="+79" swimtime="00:00:34.38" resultid="42831" heatid="45038" lane="1" entrytime="00:00:34.55" entrycourse="LCM" />
                <RESULT eventid="2682" points="299" reactiontime="+87" swimtime="00:00:39.69" resultid="42832" heatid="44895" lane="6" entrytime="00:00:39.32" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Regina Fernanda" lastname="Azevedo" birthdate="1959-11-28" gender="F" nation="POR" license="204136" swrid="5126808" athleteid="42806">
              <RESULTS>
                <RESULT eventid="2203" points="216" reactiontime="+87" swimtime="00:02:17.72" resultid="42807" heatid="44880" lane="1" entrytime="00:02:20.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="142" reactiontime="+113" swimtime="00:01:12.32" resultid="42808" heatid="45097" lane="6" entrytime="00:01:09.21" entrycourse="LCM" />
                <RESULT eventid="2460" points="144" reactiontime="+124" swimtime="00:02:43.53" resultid="42809" heatid="45118" lane="2" entrytime="00:02:37.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="278" reactiontime="+104" swimtime="00:00:59.58" resultid="42810" heatid="45023" lane="5" entrytime="00:00:58.96" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valdemar Silva" lastname="Paiva" birthdate="1977-09-18" gender="M" nation="POR" license="214138" swrid="5467379" athleteid="42857">
              <RESULTS>
                <RESULT eventid="2188" points="276" reactiontime="+96" swimtime="00:00:46.81" resultid="42858" heatid="44942" lane="1" entrytime="00:00:46.85" entrycourse="LCM" />
                <RESULT eventid="2445" points="271" reactiontime="+93" swimtime="00:01:45.94" resultid="42859" heatid="44993" lane="1" entrytime="00:01:50.03">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paula Cristina" lastname="Duarte" birthdate="1965-06-02" gender="F" nation="POR" license="207732" swrid="4885556" athleteid="42823">
              <RESULTS>
                <RESULT eventid="2607" points="290" swimtime="00:00:57.07" resultid="42824" heatid="45098" lane="4" entrytime="00:00:55.01" entrycourse="LCM" />
                <RESULT eventid="2460" points="308" swimtime="00:02:05.48" resultid="42825" heatid="45119" lane="7" entrytime="00:02:03.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="176" reactiontime="+78" swimtime="00:00:52.74" resultid="42826" heatid="45066" lane="4" entrytime="00:00:52.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filipe Jose" lastname="Baptista" birthdate="1994-01-11" gender="M" nation="POR" license="107614" swrid="4319444" athleteid="42811">
              <RESULTS>
                <RESULT eventid="1058" points="500" swimtime="00:10:56.69" resultid="42812" heatid="45085" lane="5" entrytime="00:10:11.94">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.77" />
                    <SPLIT distance="200" swimtime="00:02:35.29" />
                    <SPLIT distance="300" swimtime="00:03:58.05" />
                    <SPLIT distance="400" swimtime="00:05:22.03" />
                    <SPLIT distance="500" swimtime="00:06:46.04" />
                    <SPLIT distance="600" swimtime="00:08:11.36" />
                    <SPLIT distance="700" swimtime="00:09:35.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="558" reactiontime="+70" swimtime="00:02:19.86" resultid="42813" heatid="45095" lane="1" entrytime="00:02:27.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                    <SPLIT distance="100" swimtime="00:01:05.74" />
                    <SPLIT distance="150" swimtime="00:01:42.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" status="DNS" swimtime="00:00:00.00" resultid="42814" heatid="45114" lane="1" entrytime="00:01:03.02" entrycourse="LCM" />
                <RESULT eventid="2263" points="528" reactiontime="+73" swimtime="00:05:10.40" resultid="42815" heatid="45131" lane="7" entrytime="00:05:00.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:09.45" />
                    <SPLIT distance="150" swimtime="00:01:47.94" />
                    <SPLIT distance="200" swimtime="00:02:27.46" />
                    <SPLIT distance="250" swimtime="00:03:08.21" />
                    <SPLIT distance="300" swimtime="00:03:49.20" />
                    <SPLIT distance="350" swimtime="00:04:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="557" reactiontime="+74" swimtime="00:00:28.13" resultid="42816" heatid="45045" lane="8" entrytime="00:00:28.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Paulo" lastname="Capitao" birthdate="1996-01-31" gender="M" nation="POR" license="109592" swrid="4351797" athleteid="42817">
              <RESULTS>
                <RESULT eventid="2682" points="783" reactiontime="+73" swimtime="00:00:27.19" resultid="42818" heatid="44901" lane="2" entrytime="00:00:27.90" />
                <RESULT eventid="2323" points="622" reactiontime="+83" swimtime="00:01:06.61" resultid="42819" heatid="44930" lane="1" entrytime="00:01:04.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="694" reactiontime="+78" swimtime="00:00:58.38" resultid="42820" heatid="45115" lane="4" entrytime="00:00:58.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="527" reactiontime="+82" swimtime="00:02:35.88" resultid="42821" heatid="44982" lane="6" entrytime="00:02:31.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.56" />
                    <SPLIT distance="100" swimtime="00:01:13.83" />
                    <SPLIT distance="150" swimtime="00:01:59.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="726" reactiontime="+74" swimtime="00:00:25.75" resultid="42822" heatid="45048" lane="1" entrytime="00:00:26.06" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joana Filipa" lastname="Lamas" birthdate="1992-04-26" gender="F" nation="POR" license="13368" swrid="4074072" athleteid="42846">
              <RESULTS>
                <RESULT eventid="2607" points="528" reactiontime="+83" swimtime="00:00:40.39" resultid="42847" heatid="45103" lane="7" entrytime="00:00:40.55" entrycourse="LCM" />
                <RESULT eventid="2460" points="503" reactiontime="+82" swimtime="00:01:30.97" resultid="42848" heatid="45123" lane="1" entrytime="00:01:31.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Liza" lastname="Orioli" birthdate="1979-06-25" gender="F" nation="FRA" license="211175" swrid="5418280" athleteid="42849">
              <RESULTS>
                <RESULT eventid="2607" points="384" reactiontime="+88" swimtime="00:00:48.11" resultid="42850" heatid="45100" lane="4" entrytime="00:00:48.84" />
                <RESULT eventid="2637" points="290" reactiontime="+95" swimtime="00:01:31.11" resultid="42851" heatid="44954" lane="8" entrytime="00:01:36.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="295" reactiontime="+84" swimtime="00:00:47.56" resultid="42852" heatid="45025" lane="1" entrytime="00:00:46.74" entrycourse="LCM" />
                <RESULT eventid="2430" points="393" reactiontime="+87" swimtime="00:00:37.47" resultid="42853" heatid="45069" lane="2" entrytime="00:00:38.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ruben Manuel" lastname="Almeida" birthdate="1995-08-29" gender="M" nation="POR" license="108505" swrid="4345333" athleteid="42794">
              <RESULTS>
                <RESULT eventid="2682" points="582" reactiontime="+83" swimtime="00:00:30.02" resultid="42795" heatid="44899" lane="5" entrytime="00:00:30.27" />
                <RESULT eventid="2188" points="594" reactiontime="+79" swimtime="00:00:34.35" resultid="42796" heatid="44950" lane="2" entrytime="00:00:34.20" />
                <RESULT eventid="2415" points="618" reactiontime="+79" swimtime="00:01:00.70" resultid="42797" heatid="45114" lane="7" entrytime="00:01:02.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="456" reactiontime="+73" swimtime="00:00:34.78" resultid="42798" heatid="45020" lane="1" entrytime="00:00:35.30" />
                <RESULT eventid="2652" points="567" reactiontime="+79" swimtime="00:00:27.97" resultid="42799" heatid="45045" lane="7" entrytime="00:00:28.30" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Claudia Generosa" lastname="Gomes" birthdate="1975-10-03" gender="F" nation="POR" license="206949" swrid="5158746" athleteid="42838">
              <RESULTS>
                <RESULT eventid="2278" points="217" reactiontime="+98" swimtime="00:03:41.74" resultid="42839" heatid="44902" lane="5" entrytime="00:03:39.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.98" />
                    <SPLIT distance="100" swimtime="00:01:38.44" />
                    <SPLIT distance="150" swimtime="00:02:38.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="309" reactiontime="+102" swimtime="00:00:53.53" resultid="42840" heatid="45099" lane="2" entrytime="00:00:52.46" entrycourse="LCM" />
                <RESULT eventid="2637" points="269" reactiontime="+102" swimtime="00:01:32.79" resultid="42841" heatid="44953" lane="6" entrytime="00:01:42.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="282" reactiontime="+86" swimtime="00:02:02.05" resultid="42842" heatid="45119" lane="4" entrytime="00:01:56.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Vitor" lastname="Ferreira" birthdate="1996-05-07" gender="M" nation="POR" license="112744" swrid="4433928" athleteid="42833">
              <RESULTS>
                <RESULT eventid="2682" points="691" reactiontime="+72" swimtime="00:00:28.35" resultid="42834" heatid="44901" lane="7" entrytime="00:00:28.14" />
                <RESULT eventid="2415" points="576" reactiontime="+69" swimtime="00:01:02.14" resultid="42835" heatid="45113" lane="7" entrytime="00:01:04.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="511" reactiontime="+101" swimtime="00:00:33.48" resultid="42836" heatid="45021" lane="8" entrytime="00:00:33.40" />
                <RESULT eventid="2652" points="611" reactiontime="+73" swimtime="00:00:27.28" resultid="42837" heatid="45046" lane="4" entrytime="00:00:27.15" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique Silva" lastname="Paiva" birthdate="1967-04-08" gender="M" nation="POR" license="207623" swrid="5048945" athleteid="42854">
              <RESULTS>
                <RESULT eventid="2622" status="DNS" swimtime="00:00:00.00" resultid="42855" heatid="44873" lane="5" entrytime="00:04:22.97" entrycourse="LCM" />
                <RESULT eventid="2507" status="DNS" swimtime="00:00:00.00" resultid="42856" heatid="45090" lane="3" entrytime="00:03:58.04" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="INDANP" nation="POR" region="ANNP" clubid="41637" swrid="73274" name="Individual ANNP">
          <ATHLETES>
            <ATHLETE firstname="Alexandra Maria" lastname="Jorge" birthdate="1976-07-31" gender="F" nation="POR" license="131907" swrid="5032038" athleteid="41988">
              <RESULTS>
                <RESULT eventid="2607" points="454" reactiontime="+88" swimtime="00:00:47.10" resultid="41989" heatid="45101" lane="1" entrytime="00:00:46.98" entrycourse="LCM" />
                <RESULT eventid="2522" points="329" reactiontime="+78" swimtime="00:00:45.37" resultid="41990" heatid="45025" lane="6" entrytime="00:00:44.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Carlos" lastname="Freitas" birthdate="1963-10-24" gender="M" nation="POR" license="111877" swrid="4403503" athleteid="43609">
              <RESULTS>
                <RESULT eventid="1058" points="823" swimtime="00:10:05.03" resultid="43610" heatid="45085" lane="4" entrytime="00:09:11.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.35" />
                    <SPLIT distance="200" swimtime="00:02:27.69" />
                    <SPLIT distance="300" swimtime="00:03:43.50" />
                    <SPLIT distance="400" swimtime="00:04:59.48" />
                    <SPLIT distance="500" swimtime="00:06:16.24" />
                    <SPLIT distance="600" swimtime="00:07:33.34" />
                    <SPLIT distance="700" swimtime="00:08:50.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="861" reactiontime="+77" swimtime="00:02:16.18" resultid="43611" heatid="45096" lane="5" entrytime="00:02:07.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="100" swimtime="00:01:06.53" />
                    <SPLIT distance="150" swimtime="00:01:42.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="899" reactiontime="+79" swimtime="00:01:02.26" resultid="43612" heatid="45115" lane="5" entrytime="00:00:58.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="862" reactiontime="+79" swimtime="00:04:50.22" resultid="43613" heatid="45131" lane="5" entrytime="00:04:28.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:01:08.98" />
                    <SPLIT distance="150" swimtime="00:01:46.41" />
                    <SPLIT distance="200" swimtime="00:02:23.60" />
                    <SPLIT distance="250" swimtime="00:03:01.35" />
                    <SPLIT distance="300" swimtime="00:03:38.61" />
                    <SPLIT distance="350" swimtime="00:04:15.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rodolfo Pereira" lastname="Nunes" birthdate="1973-05-01" gender="M" nation="POR" license="25137" swrid="4575386" athleteid="41841">
              <RESULTS>
                <RESULT eventid="2537" points="609" reactiontime="+115" swimtime="00:01:12.97" resultid="41842" heatid="44888" lane="8" entrytime="00:01:16.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="664" reactiontime="+78" swimtime="00:00:30.43" resultid="41843" heatid="44899" lane="7" entrytime="00:00:30.55" entrycourse="LCM" />
                <RESULT eventid="2218" points="564" reactiontime="+83" swimtime="00:02:44.18" resultid="41844" heatid="44921" lane="7" entrytime="00:02:39.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                    <SPLIT distance="100" swimtime="00:01:21.32" />
                    <SPLIT distance="150" swimtime="00:02:03.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="687" reactiontime="+79" swimtime="00:00:33.88" resultid="41845" heatid="44950" lane="5" entrytime="00:00:32.75" entrycourse="LCM" />
                <RESULT eventid="2445" points="692" reactiontime="+87" swimtime="00:01:17.89" resultid="41846" heatid="44999" lane="3" entrytime="00:01:15.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina Santos" lastname="Silva" birthdate="1986-07-03" gender="F" nation="POR" license="23208" swrid="4064115" athleteid="41992">
              <RESULTS>
                <RESULT eventid="2203" points="650" reactiontime="+73" swimtime="00:01:20.44" resultid="41993" heatid="44883" lane="5" entrytime="00:01:10.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2552" points="607" reactiontime="+69" swimtime="00:01:18.56" resultid="41994" heatid="44924" lane="5" entrytime="00:01:06.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="628" reactiontime="+65" swimtime="00:05:28.20" resultid="41995" heatid="45013" lane="4" entrytime="00:04:53.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                    <SPLIT distance="100" swimtime="00:01:19.57" />
                    <SPLIT distance="150" swimtime="00:02:00.99" />
                    <SPLIT distance="200" swimtime="00:02:42.58" />
                    <SPLIT distance="250" swimtime="00:03:24.29" />
                    <SPLIT distance="300" swimtime="00:04:05.84" />
                    <SPLIT distance="350" swimtime="00:04:47.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="589" reactiontime="+65" swimtime="00:00:38.23" resultid="41996" heatid="45027" lane="4" entrytime="00:00:33.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ADP" nation="POR" region="ANNP" clubid="43093" swrid="66437" name="Associacao Desportiva de Penafiel" shortname="Penafiel">
          <ATHLETES>
            <ATHLETE firstname="Helder Tomas" lastname="Rocha" birthdate="1986-08-05" gender="M" nation="POR" license="203931" swrid="4235599" athleteid="44850">
              <RESULTS>
                <RESULT eventid="2652" swimtime="00:00:00.00" resultid="44851" entrytime="00:00:37.14" entrycourse="LCM" />
                <RESULT eventid="2323" points="170" reactiontime="+86" swimtime="00:01:44.92" resultid="44852" heatid="44926" lane="3" entrytime="00:01:32.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="237" reactiontime="+85" swimtime="00:01:23.88" resultid="44853" heatid="45107" lane="1" entrytime="00:01:23.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="229" reactiontime="+83" swimtime="00:03:35.82" resultid="44854" heatid="44977" lane="2" entrytime="00:03:32.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.94" />
                    <SPLIT distance="100" swimtime="00:01:41.08" />
                    <SPLIT distance="150" swimtime="00:02:48.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="237" reactiontime="+67" swimtime="00:00:43.56" resultid="44855" heatid="45017" lane="6" entrytime="00:00:45.41" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo Ricardo" lastname="Moreira" birthdate="1983-04-02" gender="M" nation="POR" license="208404" swrid="5326866" athleteid="43142">
              <RESULTS>
                <RESULT eventid="2188" status="DNS" swimtime="00:00:00.00" resultid="43143" heatid="44944" lane="8" entrytime="00:00:44.46" entrycourse="LCM" />
                <RESULT eventid="2415" status="DNS" swimtime="00:00:00.00" resultid="43144" heatid="45106" lane="7" entrytime="00:01:27.89" />
                <RESULT eventid="2445" status="DNS" swimtime="00:00:00.00" resultid="43145" heatid="44994" lane="8" entrytime="00:01:44.26" entrycourse="LCM" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="43146" heatid="45036" lane="3" entrytime="00:00:37.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel Paulo" lastname="Silva" birthdate="1971-05-03" gender="M" nation="POR" license="207402" swrid="4005722" athleteid="43156">
              <RESULTS>
                <RESULT eventid="2188" points="274" reactiontime="+100" swimtime="00:00:47.90" resultid="43157" heatid="44943" lane="7" entrytime="00:00:45.04" entrycourse="LCM" />
                <RESULT eventid="2415" points="189" reactiontime="+97" swimtime="00:01:38.92" resultid="43158" heatid="45105" lane="5" entrytime="00:01:30.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.59" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="720 - Toque alternado na viragem aos 50 m - SW 7.6" eventid="2445" reactiontime="+93" status="DSQ" swimtime="00:01:55.56" resultid="43159" heatid="44994" lane="6" entrytime="00:01:43.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="199" reactiontime="+88" swimtime="00:00:43.00" resultid="43160" heatid="45034" lane="2" entrytime="00:00:43.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Manuel" lastname="Ventura" birthdate="1983-12-24" gender="M" nation="POR" license="153165" swrid="5113030" athleteid="43166">
              <RESULTS>
                <RESULT eventid="2188" points="376" reactiontime="+115" swimtime="00:00:40.46" resultid="43167" heatid="44942" lane="5" entrytime="00:00:45.54" />
                <RESULT eventid="2415" points="354" reactiontime="+94" swimtime="00:01:13.43" resultid="43168" heatid="45109" lane="1" entrytime="00:01:16.26">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="355" reactiontime="+99" swimtime="00:01:33.81" resultid="43169" heatid="44995" lane="3" entrytime="00:01:37.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" status="DNS" swimtime="00:00:00.00" resultid="43170" heatid="45126" lane="2" entrytime="00:07:15.45" entrycourse="LCM" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="43171" heatid="45037" lane="6" entrytime="00:00:35.69" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabio Andre" lastname="Madureira" birthdate="1990-05-19" gender="M" nation="POR" license="15910" swrid="4073863" athleteid="43133">
              <RESULTS>
                <RESULT eventid="2188" points="554" reactiontime="+84" swimtime="00:00:35.05" resultid="43134" heatid="44950" lane="6" entrytime="00:00:33.89" entrycourse="LCM" />
                <RESULT eventid="2385" points="462" reactiontime="+85" swimtime="00:02:50.20" resultid="43135" heatid="44979" lane="7" entrytime="00:03:00.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                    <SPLIT distance="100" swimtime="00:01:24.93" />
                    <SPLIT distance="150" swimtime="00:02:11.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="358" reactiontime="+89" swimtime="00:05:49.82" resultid="43136" heatid="45129" lane="1" entrytime="00:05:53.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                    <SPLIT distance="100" swimtime="00:01:20.10" />
                    <SPLIT distance="150" swimtime="00:02:04.82" />
                    <SPLIT distance="200" swimtime="00:02:50.31" />
                    <SPLIT distance="250" swimtime="00:03:35.21" />
                    <SPLIT distance="300" swimtime="00:04:22.17" />
                    <SPLIT distance="350" swimtime="00:05:09.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" points="343" reactiontime="+88" swimtime="00:03:09.03" resultid="43137" heatid="45029" lane="3" entrytime="00:03:20.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.91" />
                    <SPLIT distance="100" swimtime="00:01:34.54" />
                    <SPLIT distance="150" swimtime="00:02:20.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Maria" lastname="Ramalho" birthdate="1952-09-01" gender="M" nation="POR" license="211689" swrid="5377395" athleteid="43152">
              <RESULTS>
                <RESULT eventid="2188" points="223" reactiontime="+125" swimtime="00:00:56.87" resultid="43153" heatid="44939" lane="2" entrytime="00:00:57.86" entrycourse="LCM" />
                <RESULT eventid="2445" points="242" reactiontime="+117" swimtime="00:02:12.10" resultid="43154" heatid="44990" lane="4" entrytime="00:02:17.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="141" reactiontime="+122" swimtime="00:00:54.52" resultid="43155" heatid="45033" lane="7" entrytime="00:01:00.56" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Joaquim" lastname="Moreira" birthdate="1987-06-05" gender="M" nation="POR" license="131844" swrid="5041332" athleteid="43147">
              <RESULTS>
                <RESULT eventid="2323" points="323" reactiontime="+78" swimtime="00:01:22.61" resultid="43148" heatid="44928" lane="8" entrytime="00:01:14.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="454" reactiontime="+68" swimtime="00:01:06.11" resultid="43149" heatid="45113" lane="8" entrytime="00:01:04.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="403 - Falsa partida - SW 4.4" eventid="2385" reactiontime="+78" status="DSQ" swimtime="00:02:57.05" resultid="43150" heatid="44981" lane="7" entrytime="00:02:45.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                    <SPLIT distance="100" swimtime="00:01:23.92" />
                    <SPLIT distance="150" swimtime="00:02:14.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="347" reactiontime="+88" swimtime="00:01:30.91" resultid="43151" heatid="44998" lane="1" entrytime="00:01:24.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jaime Antonio" lastname="Soares" birthdate="1987-07-02" gender="M" nation="POR" license="208104" swrid="5320572" athleteid="43161">
              <RESULTS>
                <RESULT eventid="2188" points="253" reactiontime="+107" swimtime="00:00:45.48" resultid="43162" heatid="44942" lane="6" entrytime="00:00:46.05" entrycourse="LCM" />
                <RESULT eventid="2415" points="333" reactiontime="+97" swimtime="00:01:13.29" resultid="43163" heatid="45108" lane="4" entrytime="00:01:17.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="270" reactiontime="+109" swimtime="00:00:40.22" resultid="43164" heatid="45017" lane="5" entrytime="00:00:44.87" />
                <RESULT eventid="2652" points="341" reactiontime="+96" swimtime="00:00:33.26" resultid="43165" heatid="45038" lane="8" entrytime="00:00:34.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Vieira" lastname="Moreira" birthdate="1957-09-29" gender="F" nation="POR" license="205072" swrid="5229971" athleteid="43138">
              <RESULTS>
                <RESULT eventid="2637" points="108" swimtime="00:02:27.21" resultid="43139" heatid="44951" lane="4" entrytime="00:02:16.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="133" reactiontime="+91" swimtime="00:01:16.21" resultid="43140" heatid="45023" lane="7" entrytime="00:01:12.75" entrycourse="LCM" />
                <RESULT eventid="2430" points="131" swimtime="00:01:01.28" resultid="43141" heatid="45065" lane="4" entrytime="00:01:05.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LSC" nation="POR" region="ANNP" clubid="41929" swrid="65800" name="Leixoes Sport Club" shortname="Leixoes">
          <ATHLETES>
            <ATHLETE firstname="Luis Filipe" lastname="Rato" birthdate="1981-01-05" gender="M" nation="POR" license="26260" swrid="4074138" athleteid="43941">
              <RESULTS>
                <RESULT eventid="2537" points="483" reactiontime="+72" swimtime="00:01:18.23" resultid="43942" heatid="44887" lane="5" entrytime="00:01:19.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="515" reactiontime="+82" swimtime="00:02:45.16" resultid="43943" heatid="44980" lane="7" entrytime="00:02:54.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:18.00" />
                    <SPLIT distance="150" swimtime="00:02:06.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernando Santos" lastname="Moreira" birthdate="1994-09-03" gender="M" nation="POR" license="15824" swrid="4561322" athleteid="43932">
              <RESULTS>
                <RESULT eventid="2682" points="704" reactiontime="+85" swimtime="00:00:28.18" resultid="43933" heatid="44900" lane="4" entrytime="00:00:28.61" entrycourse="LCM" />
                <RESULT eventid="2323" points="654" reactiontime="+81" swimtime="00:01:05.49" resultid="43934" heatid="44929" lane="6" entrytime="00:01:06.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="651" reactiontime="+81" swimtime="00:00:59.65" resultid="43935" heatid="45115" lane="6" entrytime="00:00:59.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="659" reactiontime="+81" swimtime="00:00:26.60" resultid="43936" heatid="45048" lane="8" entrytime="00:00:26.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Miguel" lastname="Antunes" birthdate="1968-03-18" gender="M" nation="POR" license="206896" swrid="5276395" athleteid="43830">
              <RESULTS>
                <RESULT eventid="2537" points="196" reactiontime="+72" swimtime="00:01:53.19" resultid="43831" heatid="44885" lane="2" entrytime="00:01:55.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="231" reactiontime="+116" swimtime="00:03:27.25" resultid="43832" heatid="45091" lane="7" entrytime="00:03:29.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.95" />
                    <SPLIT distance="100" swimtime="00:01:39.39" />
                    <SPLIT distance="150" swimtime="00:02:35.91" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="603 - Após viragem saiu em posição ventral aos 100 m - SW 6.2" eventid="2218" reactiontime="+83" status="DSQ" swimtime="00:04:07.90" resultid="43833" heatid="44917" lane="7" entrytime="00:04:23.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.03" />
                    <SPLIT distance="100" swimtime="00:02:04.45" />
                    <SPLIT distance="150" swimtime="00:03:10.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="254" reactiontime="+117" swimtime="00:01:29.78" resultid="43834" heatid="45105" lane="6" entrytime="00:01:32.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="229" reactiontime="+126" swimtime="00:07:16.59" resultid="43835" heatid="45125" lane="5" entrytime="00:07:45.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.31" />
                    <SPLIT distance="100" swimtime="00:01:43.90" />
                    <SPLIT distance="150" swimtime="00:02:39.56" />
                    <SPLIT distance="200" swimtime="00:03:36.28" />
                    <SPLIT distance="250" swimtime="00:04:32.84" />
                    <SPLIT distance="300" swimtime="00:05:29.11" />
                    <SPLIT distance="350" swimtime="00:06:24.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Bruno" lastname="Meneses" birthdate="1962-11-29" gender="M" nation="POR" license="132358" swrid="5065803" athleteid="43922">
              <RESULTS>
                <RESULT eventid="2537" status="DNS" swimtime="00:00:00.00" resultid="43923" heatid="44886" lane="5" entrytime="00:01:33.16" entrycourse="LCM" />
                <RESULT eventid="2682" status="DNS" swimtime="00:00:00.00" resultid="43924" heatid="44895" lane="4" entrytime="00:00:37.72" entrycourse="LCM" />
                <RESULT eventid="2415" status="DNS" swimtime="00:00:00.00" resultid="43925" heatid="45110" lane="3" entrytime="00:01:11.06" entrycourse="LCM" />
                <RESULT eventid="2293" points="396" reactiontime="+70" swimtime="00:00:42.63" resultid="43926" heatid="45018" lane="1" entrytime="00:00:43.03" entrycourse="LCM" />
                <RESULT eventid="2652" points="548" reactiontime="+103" swimtime="00:00:32.51" resultid="43927" heatid="45040" lane="5" entrytime="00:00:31.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Manuel" lastname="Fonseca" birthdate="1987-07-18" gender="M" nation="POR" license="25159" swrid="4064552" athleteid="43891">
              <RESULTS>
                <RESULT eventid="2323" points="523" reactiontime="+82" swimtime="00:01:10.33" resultid="43892" heatid="44929" lane="5" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="575" reactiontime="+81" swimtime="00:02:38.21" resultid="43893" heatid="44982" lane="7" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.55" />
                    <SPLIT distance="100" swimtime="00:01:13.12" />
                    <SPLIT distance="150" swimtime="00:01:59.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="601" reactiontime="+80" swimtime="00:00:27.55" resultid="43894" heatid="45044" lane="4" entrytime="00:00:28.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Graca Maria" lastname="Almeida" birthdate="1973-08-18" gender="F" nation="POR" license="124702" swrid="4004774" athleteid="43827">
              <RESULTS>
                <RESULT eventid="2308" status="WDR" swimtime="00:00:00.00" resultid="43828" entrytime="00:03:13.43" entrycourse="LCM" />
                <RESULT eventid="2522" points="402" reactiontime="+89" swimtime="00:00:42.44" resultid="43829" heatid="45025" lane="5" entrytime="00:00:41.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Antonio" lastname="Ferreira" birthdate="1958-07-17" gender="M" nation="POR" license="214085" swrid="5465976" athleteid="43879">
              <RESULTS>
                <RESULT eventid="1058" points="295" swimtime="00:15:39.86" resultid="43880" heatid="45080" lane="3" entrytime="00:16:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.78" />
                    <SPLIT distance="200" swimtime="00:03:48.74" />
                    <SPLIT distance="300" swimtime="00:05:48.18" />
                    <SPLIT distance="400" swimtime="00:07:46.89" />
                    <SPLIT distance="500" swimtime="00:09:45.40" />
                    <SPLIT distance="600" swimtime="00:11:46.04" />
                    <SPLIT distance="700" swimtime="00:13:45.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="146" reactiontime="+106" swimtime="00:00:55.27" resultid="43881" heatid="44893" lane="7" entrytime="00:00:55.00" />
                <RESULT eventid="2218" points="250" reactiontime="+98" swimtime="00:04:18.61" resultid="43882" heatid="44917" lane="2" entrytime="00:04:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.24" />
                    <SPLIT distance="100" swimtime="00:02:06.90" />
                    <SPLIT distance="150" swimtime="00:03:13.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="310" reactiontime="+116" swimtime="00:07:22.67" resultid="43883" heatid="45126" lane="7" entrytime="00:07:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.14" />
                    <SPLIT distance="100" swimtime="00:01:39.30" />
                    <SPLIT distance="150" swimtime="00:02:35.81" />
                    <SPLIT distance="200" swimtime="00:03:32.75" />
                    <SPLIT distance="250" swimtime="00:04:30.60" />
                    <SPLIT distance="300" swimtime="00:05:29.77" />
                    <SPLIT distance="350" swimtime="00:06:29.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="299" reactiontime="+101" swimtime="00:01:55.07" resultid="43884" heatid="44991" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Pedro" lastname="Castro" birthdate="1974-06-10" gender="M" nation="POR" license="132355" swrid="5065798" athleteid="43853">
              <RESULTS>
                <RESULT eventid="2682" status="DNS" swimtime="00:00:00.00" resultid="43854" heatid="44896" lane="8" entrytime="00:00:37.28" entrycourse="LCM" />
                <RESULT eventid="2415" status="DNS" swimtime="00:00:00.00" resultid="43855" heatid="45110" lane="1" entrytime="00:01:12.24" entrycourse="LCM" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="43856" heatid="45040" lane="4" entrytime="00:00:31.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo Amorim" lastname="Rego" birthdate="1984-06-24" gender="M" nation="POR" license="15954" swrid="4064560" athleteid="43944">
              <RESULTS>
                <RESULT eventid="2218" points="613" reactiontime="+85" swimtime="00:02:36.75" resultid="43945" heatid="44921" lane="3" entrytime="00:02:29.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="100" swimtime="00:01:13.23" />
                    <SPLIT distance="150" swimtime="00:01:53.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="714" reactiontime="+84" swimtime="00:02:27.77" resultid="43946" heatid="44982" lane="5" entrytime="00:02:23.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.74" />
                    <SPLIT distance="100" swimtime="00:01:08.92" />
                    <SPLIT distance="150" swimtime="00:01:50.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="590" reactiontime="+95" swimtime="00:00:32.18" resultid="43947" heatid="45022" lane="3" entrytime="00:00:31.05" entrycourse="LCM" />
                <RESULT eventid="2445" points="662" reactiontime="+82" swimtime="00:01:16.24" resultid="43948" heatid="44999" lane="5" entrytime="00:01:13.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="667" reactiontime="+79" swimtime="00:05:26.11" resultid="43949" heatid="45062" lane="5" entrytime="00:05:06.20">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                    <SPLIT distance="100" swimtime="00:01:12.19" />
                    <SPLIT distance="150" swimtime="00:01:55.22" />
                    <SPLIT distance="200" swimtime="00:02:38.56" />
                    <SPLIT distance="250" swimtime="00:03:22.42" />
                    <SPLIT distance="300" swimtime="00:04:07.71" />
                    <SPLIT distance="350" swimtime="00:04:47.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Luisa" lastname="Garcia" birthdate="1970-10-05" gender="F" nation="POR" license="214120" swrid="5465977" athleteid="43898">
              <RESULTS>
                <RESULT eventid="1060" points="190" swimtime="00:17:09.05" resultid="43899" heatid="45074" lane="3" entrytime="00:18:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:04.07" />
                    <SPLIT distance="200" swimtime="00:04:10.23" />
                    <SPLIT distance="300" swimtime="00:06:17.18" />
                    <SPLIT distance="400" swimtime="00:08:25.66" />
                    <SPLIT distance="500" swimtime="00:10:34.36" />
                    <SPLIT distance="600" swimtime="00:12:43.01" />
                    <SPLIT distance="700" swimtime="00:14:56.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2173" points="384" swimtime="00:04:11.94" resultid="43900" heatid="45087" lane="2" entrytime="00:04:25.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.36" />
                    <SPLIT distance="100" swimtime="00:02:02.27" />
                    <SPLIT distance="150" swimtime="00:03:06.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" status="DNS" swimtime="00:00:00.00" resultid="43901" heatid="45099" lane="8" entrytime="00:00:54.59" entrycourse="LCM" />
                <RESULT eventid="2637" points="174" reactiontime="+115" swimtime="00:01:53.29" resultid="43902" heatid="44952" lane="5" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Carmo" lastname="Rocha" birthdate="1954-08-19" gender="F" nation="POR" license="118886" swrid="4590378" athleteid="43953">
              <RESULTS>
                <RESULT eventid="2173" status="DNS" swimtime="00:00:00.00" resultid="43954" heatid="45086" lane="3" entrytime="00:05:02.41" entrycourse="LCM" />
                <RESULT eventid="2607" status="DNS" swimtime="00:00:00.00" resultid="43955" heatid="45097" lane="5" entrytime="00:01:05.42" entrycourse="LCM" />
                <RESULT eventid="2522" points="84" reactiontime="+93" swimtime="00:01:32.50" resultid="43956" heatid="45023" lane="1" entrytime="00:01:35.50" entrycourse="LCM" />
                <RESULT eventid="2460" status="DNS" swimtime="00:00:00.00" resultid="43957" heatid="45118" lane="6" entrytime="00:02:27.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hugo Rafael" lastname="Guedes" birthdate="1976-10-22" gender="M" nation="POR" license="204930" swrid="5220479" athleteid="43909">
              <RESULTS>
                <RESULT eventid="2188" points="342" reactiontime="+88" swimtime="00:00:42.72" resultid="43910" heatid="44945" lane="5" entrytime="00:00:41.93" entrycourse="LCM" />
                <RESULT eventid="2415" points="279" reactiontime="+92" swimtime="00:01:25.47" resultid="43911" heatid="45106" lane="3" entrytime="00:01:26.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="317" reactiontime="+96" swimtime="00:01:40.98" resultid="43912" heatid="44995" lane="7" entrytime="00:01:39.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="338" reactiontime="+83" swimtime="00:00:35.69" resultid="43913" heatid="45035" lane="1" entrytime="00:00:41.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joana Maria" lastname="Faria" birthdate="1974-06-08" gender="F" nation="POR" license="128933" swrid="4940519" athleteid="43868">
              <RESULTS>
                <RESULT eventid="2607" points="603" reactiontime="+97" swimtime="00:00:42.85" resultid="43869" heatid="45102" lane="5" entrytime="00:00:42.15" entrycourse="LCM" />
                <RESULT eventid="2233" points="511" reactiontime="+102" swimtime="00:03:10.09" resultid="43870" heatid="44974" lane="1" entrytime="00:03:02.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                    <SPLIT distance="100" swimtime="00:01:30.01" />
                    <SPLIT distance="150" swimtime="00:02:23.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2667" points="422" reactiontime="+98" swimtime="00:03:27.61" resultid="43871" heatid="45031" lane="5" entrytime="00:03:23.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                    <SPLIT distance="100" swimtime="00:01:37.61" />
                    <SPLIT distance="150" swimtime="00:02:32.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="594" reactiontime="+95" swimtime="00:01:35.26" resultid="43872" heatid="45123" lane="8" entrytime="00:01:32.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="540" reactiontime="+94" swimtime="00:00:34.09" resultid="43873" heatid="45071" lane="6" entrytime="00:00:33.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno Daniel" lastname="Monteiro" birthdate="1988-06-19" gender="M" nation="POR" license="26069" swrid="4064548" athleteid="43928">
              <RESULTS>
                <RESULT eventid="2622" points="748" reactiontime="+75" swimtime="00:02:38.01" resultid="43929" heatid="44879" lane="4" entrytime="00:02:38.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:17.21" />
                    <SPLIT distance="150" swimtime="00:01:59.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="801" reactiontime="+77" swimtime="00:00:30.99" resultid="43930" heatid="44950" lane="4" entrytime="00:00:30.67" entrycourse="LCM" />
                <RESULT eventid="2445" points="797" reactiontime="+73" swimtime="00:01:08.92" resultid="43931" heatid="44999" lane="4" entrytime="00:01:08.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nuno Alexandre" lastname="Viseu" birthdate="1977-12-14" gender="M" nation="POR" license="205761" swrid="5260691" athleteid="43978">
              <RESULTS>
                <RESULT eventid="2188" points="287" reactiontime="+99" swimtime="00:00:46.25" resultid="43979" heatid="44942" lane="2" entrytime="00:00:46.28" entrycourse="LCM" />
                <RESULT eventid="2385" points="195" reactiontime="+99" swimtime="00:03:48.25" resultid="43980" heatid="44976" lane="6" entrytime="00:03:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.21" />
                    <SPLIT distance="100" swimtime="00:01:54.95" />
                    <SPLIT distance="150" swimtime="00:02:57.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="146" reactiontime="+74" swimtime="00:00:53.85" resultid="43981" heatid="45015" lane="7" entrytime="00:00:56.49" entrycourse="LCM" />
                <RESULT eventid="2652" points="392" reactiontime="+100" swimtime="00:00:33.58" resultid="43982" heatid="45039" lane="1" entrytime="00:00:33.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edgar Francisco" lastname="Ribeiro" birthdate="1991-08-02" gender="M" nation="POR" license="208133" swrid="5411288" athleteid="43950">
              <RESULTS>
                <RESULT eventid="1058" points="253" swimtime="00:12:51.86" resultid="43951" heatid="45083" lane="1" entrytime="00:12:48.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.92" />
                    <SPLIT distance="200" swimtime="00:03:02.66" />
                    <SPLIT distance="300" swimtime="00:04:40.14" />
                    <SPLIT distance="400" swimtime="00:06:18.76" />
                    <SPLIT distance="500" swimtime="00:07:58.89" />
                    <SPLIT distance="600" swimtime="00:09:37.94" />
                    <SPLIT distance="700" swimtime="00:11:16.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" status="DNS" swimtime="00:00:00.00" resultid="43952" heatid="44895" lane="3" entrytime="00:00:39.22" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Manuel" lastname="Baptista" birthdate="1969-09-20" gender="M" nation="POR" license="130027" swrid="4989261" athleteid="43836">
              <RESULTS>
                <RESULT eventid="2622" points="333" reactiontime="+117" swimtime="00:03:50.90" resultid="43837" heatid="44875" lane="1" entrytime="00:03:45.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.36" />
                    <SPLIT distance="100" swimtime="00:01:51.47" />
                    <SPLIT distance="150" swimtime="00:02:52.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2323" points="119" reactiontime="+132" swimtime="00:02:09.46" resultid="43838" heatid="44925" lane="2" entrytime="00:02:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="188" reactiontime="+129" swimtime="00:04:11.43" resultid="43839" heatid="44975" lane="4" entrytime="00:04:09.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.43" />
                    <SPLIT distance="100" swimtime="00:02:16.08" />
                    <SPLIT distance="150" swimtime="00:03:14.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="308" reactiontime="+126" swimtime="00:01:47.34" resultid="43840" heatid="44994" lane="7" entrytime="00:01:43.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="203" reactiontime="+126" swimtime="00:08:59.52" resultid="43841" heatid="45059" lane="7" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.23" />
                    <SPLIT distance="100" swimtime="00:02:11.37" />
                    <SPLIT distance="150" swimtime="00:03:33.71" />
                    <SPLIT distance="200" swimtime="00:04:58.17" />
                    <SPLIT distance="250" swimtime="00:05:57.97" />
                    <SPLIT distance="300" swimtime="00:07:01.20" />
                    <SPLIT distance="350" swimtime="00:08:01.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel Jose" lastname="Ferreira" birthdate="1970-07-27" gender="M" nation="POR" license="119657" swrid="4607066" athleteid="43885">
              <RESULTS>
                <RESULT eventid="2218" points="445" reactiontime="+79" swimtime="00:03:14.18" resultid="43886" heatid="44920" lane="8" entrytime="00:03:07.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                    <SPLIT distance="100" swimtime="00:01:33.59" />
                    <SPLIT distance="150" swimtime="00:02:25.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="528" reactiontime="+84" swimtime="00:01:10.31" resultid="43887" heatid="45111" lane="5" entrytime="00:01:07.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="380" reactiontime="+82" swimtime="00:03:19.04" resultid="43888" heatid="44977" lane="3" entrytime="00:03:22.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                    <SPLIT distance="100" swimtime="00:01:35.26" />
                    <SPLIT distance="150" swimtime="00:02:37.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="489" reactiontime="+74" swimtime="00:00:37.77" resultid="43889" heatid="45019" lane="3" entrytime="00:00:37.42" entrycourse="LCM" />
                <RESULT eventid="2652" points="568" reactiontime="+76" swimtime="00:00:30.33" resultid="43890" heatid="45042" lane="2" entrytime="00:00:30.11" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre Filipe" lastname="Couto" birthdate="1991-04-07" gender="M" nation="POR" license="23958" swrid="4269384" athleteid="43857">
              <RESULTS>
                <RESULT eventid="2682" status="DNS" swimtime="00:00:00.00" resultid="43858" heatid="44899" lane="1" entrytime="00:00:30.72" entrycourse="LCM" />
                <RESULT eventid="2507" status="DNS" swimtime="00:00:00.00" resultid="43859" heatid="45093" lane="8" entrytime="00:02:50.95" entrycourse="LCM" />
                <RESULT eventid="2415" status="DNS" swimtime="00:00:00.00" resultid="43860" heatid="45114" lane="5" entrytime="00:01:01.14" entrycourse="LCM" />
                <RESULT eventid="2263" status="DNS" swimtime="00:00:00.00" resultid="43861" heatid="45129" lane="7" entrytime="00:05:51.53" entrycourse="LCM" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="43862" heatid="45043" lane="4" entrytime="00:00:28.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Santos" lastname="Fernandes" birthdate="1962-03-28" gender="F" nation="POR" license="105263" swrid="4246947" athleteid="43874">
              <RESULTS>
                <RESULT eventid="1060" points="325" swimtime="00:14:39.53" resultid="43875" heatid="45077" lane="8" entrytime="00:14:17.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.48" />
                    <SPLIT distance="200" swimtime="00:03:31.71" />
                    <SPLIT distance="300" swimtime="00:05:22.92" />
                    <SPLIT distance="400" swimtime="00:07:15.55" />
                    <SPLIT distance="500" swimtime="00:09:07.49" />
                    <SPLIT distance="600" swimtime="00:10:59.85" />
                    <SPLIT distance="700" swimtime="00:12:50.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2173" points="491" swimtime="00:03:59.95" resultid="43876" heatid="45088" lane="3" entrytime="00:03:50.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.44" />
                    <SPLIT distance="100" swimtime="00:01:56.90" />
                    <SPLIT distance="150" swimtime="00:02:57.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="333" reactiontime="+108" swimtime="00:06:59.38" resultid="43877" heatid="45011" lane="8" entrytime="00:06:57.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.03" />
                    <SPLIT distance="100" swimtime="00:01:38.16" />
                    <SPLIT distance="150" swimtime="00:02:31.56" />
                    <SPLIT distance="200" swimtime="00:03:25.60" />
                    <SPLIT distance="250" swimtime="00:04:19.61" />
                    <SPLIT distance="300" swimtime="00:05:13.63" />
                    <SPLIT distance="350" swimtime="00:06:07.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="452" reactiontime="+107" swimtime="00:01:50.39" resultid="43878" heatid="45121" lane="7" entrytime="00:01:46.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Adriana" lastname="Viseu" birthdate="1966-03-13" gender="F" nation="POR" license="26830" swrid="4576017" athleteid="43972">
              <RESULTS>
                <RESULT eventid="2607" points="535" reactiontime="+83" swimtime="00:00:46.56" resultid="43973" heatid="45101" lane="6" entrytime="00:00:45.51" entrycourse="LCM" />
                <RESULT eventid="2637" points="416" reactiontime="+83" swimtime="00:01:25.27" resultid="43974" heatid="44955" lane="3" entrytime="00:01:21.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="354" reactiontime="+89" swimtime="00:06:50.74" resultid="43975" heatid="45011" lane="7" entrytime="00:06:56.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.18" />
                    <SPLIT distance="100" swimtime="00:01:32.39" />
                    <SPLIT distance="150" swimtime="00:02:24.35" />
                    <SPLIT distance="200" swimtime="00:03:17.22" />
                    <SPLIT distance="250" swimtime="00:04:11.22" />
                    <SPLIT distance="300" swimtime="00:05:04.06" />
                    <SPLIT distance="350" swimtime="00:05:58.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="525" reactiontime="+93" swimtime="00:01:45.03" resultid="43976" heatid="45121" lane="3" entrytime="00:01:41.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="491" reactiontime="+85" swimtime="00:00:37.53" resultid="43977" heatid="45070" lane="8" entrytime="00:00:36.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana DAlte" lastname="Guedes" birthdate="1980-11-23" gender="F" nation="POR" license="121739" swrid="4703108" athleteid="43903">
              <RESULTS>
                <RESULT eventid="2203" points="349" reactiontime="+70" swimtime="00:01:39.48" resultid="43904" heatid="44882" lane="7" entrytime="00:01:38.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2278" points="427" reactiontime="+95" swimtime="00:02:54.75" resultid="43905" heatid="44904" lane="3" entrytime="00:02:54.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:23.44" />
                    <SPLIT distance="150" swimtime="00:02:09.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="451" reactiontime="+94" swimtime="00:01:18.62" resultid="43906" heatid="44956" lane="8" entrytime="00:01:18.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="455" reactiontime="+95" swimtime="00:06:07.53" resultid="43907" heatid="45012" lane="5" entrytime="00:06:14.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                    <SPLIT distance="100" swimtime="00:01:25.06" />
                    <SPLIT distance="150" swimtime="00:02:12.87" />
                    <SPLIT distance="200" swimtime="00:03:00.68" />
                    <SPLIT distance="250" swimtime="00:03:48.35" />
                    <SPLIT distance="300" swimtime="00:04:35.81" />
                    <SPLIT distance="350" swimtime="00:05:23.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="316" reactiontime="+78" swimtime="00:00:46.47" resultid="43908" heatid="45025" lane="2" entrytime="00:00:45.19" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joana Filipa" lastname="Rosas" birthdate="1995-01-08" gender="F" nation="POR" license="102023" swrid="4123417" athleteid="43958">
              <RESULTS>
                <RESULT eventid="1060" points="524" swimtime="00:11:25.14" resultid="43959" heatid="45078" lane="5" entrytime="00:11:14.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                    <SPLIT distance="200" swimtime="00:02:42.71" />
                    <SPLIT distance="300" swimtime="00:04:10.04" />
                    <SPLIT distance="400" swimtime="00:05:38.75" />
                    <SPLIT distance="500" swimtime="00:07:06.59" />
                    <SPLIT distance="600" swimtime="00:08:34.41" />
                    <SPLIT distance="700" swimtime="00:10:01.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="563" reactiontime="+96" swimtime="00:02:52.64" resultid="43960" heatid="44974" lane="6" entrytime="00:02:53.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                    <SPLIT distance="100" swimtime="00:01:21.65" />
                    <SPLIT distance="150" swimtime="00:02:12.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helder Ricardo" lastname="Machado" birthdate="1976-07-03" gender="M" nation="POR" license="132360" swrid="5065802" athleteid="43914">
              <RESULTS>
                <RESULT eventid="2248" points="248" reactiontime="+107" swimtime="00:08:01.10" resultid="43915" heatid="45059" lane="6" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.90" />
                    <SPLIT distance="100" swimtime="00:01:46.77" />
                    <SPLIT distance="150" swimtime="00:02:55.74" />
                    <SPLIT distance="200" swimtime="00:04:02.25" />
                    <SPLIT distance="250" swimtime="00:05:00.85" />
                    <SPLIT distance="300" swimtime="00:06:02.76" />
                    <SPLIT distance="350" swimtime="00:07:01.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Azucena" lastname="Canora Marin" birthdate="1960-03-14" gender="F" nation="ESP" license="214254" swrid="5236524" athleteid="43847">
              <RESULTS>
                <RESULT eventid="2173" points="450" swimtime="00:04:15.29" resultid="43848" heatid="45087" lane="3" entrytime="00:04:10.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.27" />
                    <SPLIT distance="100" swimtime="00:02:00.10" />
                    <SPLIT distance="150" swimtime="00:03:07.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2338" points="281" reactiontime="+93" swimtime="00:00:50.98" resultid="43849" heatid="44890" lane="1" entrytime="00:00:50.96" entrycourse="LCM" />
                <RESULT eventid="2552" points="260" reactiontime="+84" swimtime="00:02:07.25" resultid="43850" heatid="44923" lane="6" entrytime="00:01:59.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="452" reactiontime="+78" swimtime="00:01:31.58" resultid="43851" heatid="44955" lane="1" entrytime="00:01:27.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="514" reactiontime="+90" swimtime="00:07:15.37" resultid="43852" heatid="45010" lane="7" entrytime="00:07:21.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.25" />
                    <SPLIT distance="100" swimtime="00:01:39.83" />
                    <SPLIT distance="150" swimtime="00:02:35.50" />
                    <SPLIT distance="200" swimtime="00:03:31.53" />
                    <SPLIT distance="250" swimtime="00:04:28.03" />
                    <SPLIT distance="300" swimtime="00:05:24.67" />
                    <SPLIT distance="350" swimtime="00:06:21.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Henrique" lastname="Seara" birthdate="1963-10-01" gender="M" nation="POR" license="131833" swrid="5041337" athleteid="43961">
              <RESULTS>
                <RESULT eventid="2622" points="255" reactiontime="+87" swimtime="00:04:17.72" resultid="43962" heatid="44874" lane="7" entrytime="00:04:12.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.54" />
                    <SPLIT distance="100" swimtime="00:01:56.86" />
                    <SPLIT distance="150" swimtime="00:03:05.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2537" points="155" reactiontime="+78" swimtime="00:02:06.95" resultid="43963" heatid="44885" lane="8" entrytime="00:02:05.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.98" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="403 - Falsa partida - SW 4.4" eventid="2188" reactiontime="+77" status="DSQ" swimtime="00:00:49.87" resultid="43964" heatid="44939" lane="4" entrytime="00:00:51.68" entrycourse="LCM" />
                <RESULT eventid="2293" points="167" reactiontime="+86" swimtime="00:00:56.84" resultid="43965" heatid="45016" lane="8" entrytime="00:00:53.96" entrycourse="LCM" />
                <RESULT eventid="2445" points="234" reactiontime="+105" swimtime="00:01:57.76" resultid="43966" heatid="44992" lane="2" entrytime="00:01:57.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cristina Isabel" lastname="Moura" birthdate="1963-07-31" gender="F" nation="POR" license="200762" swrid="5157468" athleteid="43937">
              <RESULTS>
                <RESULT eventid="2607" points="420" reactiontime="+98" swimtime="00:00:50.47" resultid="43938" heatid="45099" lane="6" entrytime="00:00:52.25" entrycourse="LCM" />
                <RESULT eventid="2522" points="285" reactiontime="+129" swimtime="00:00:54.28" resultid="43939" heatid="45024" lane="7" entrytime="00:00:53.83" entrycourse="LCM" />
                <RESULT eventid="2430" points="312" reactiontime="+109" swimtime="00:00:43.63" resultid="43940" heatid="45067" lane="5" entrytime="00:00:44.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Pedro" lastname="Machado" birthdate="1986-11-09" gender="M" nation="POR" license="125910" swrid="4558986" athleteid="43916">
              <RESULTS>
                <RESULT eventid="2682" points="716" reactiontime="+82" swimtime="00:00:28.52" resultid="43917" heatid="44900" lane="3" entrytime="00:00:29.08" entrycourse="LCM" />
                <RESULT eventid="2323" points="597" reactiontime="+82" swimtime="00:01:09.15" resultid="43918" heatid="44929" lane="3" entrytime="00:01:06.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="576" reactiontime="+84" swimtime="00:02:38.77" resultid="43919" heatid="44981" lane="3" entrytime="00:02:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                    <SPLIT distance="100" swimtime="00:01:11.33" />
                    <SPLIT distance="150" swimtime="00:01:59.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="575" reactiontime="+104" swimtime="00:00:32.44" resultid="43920" heatid="45021" lane="5" entrytime="00:00:33.00" />
                <RESULT eventid="2652" points="558" reactiontime="+86" swimtime="00:00:28.58" resultid="43921" heatid="45043" lane="3" entrytime="00:00:29.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elsa Maria" lastname="Fumega" birthdate="1978-08-21" gender="F" nation="POR" license="119665" swrid="4607079" athleteid="43895">
              <RESULTS>
                <RESULT eventid="2607" points="583" reactiontime="+82" swimtime="00:00:41.85" resultid="43896" heatid="45102" lane="6" entrytime="00:00:43.36" entrycourse="LCM" />
                <RESULT eventid="2233" points="485" reactiontime="+85" swimtime="00:03:12.65" resultid="43897" heatid="44973" lane="2" entrytime="00:03:12.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                    <SPLIT distance="100" swimtime="00:01:32.21" />
                    <SPLIT distance="150" swimtime="00:02:26.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raquel Alexandra" lastname="Silva" birthdate="1991-06-04" gender="F" nation="POR" license="26074" swrid="4061684" athleteid="43967">
              <RESULTS>
                <RESULT eventid="2552" points="603" reactiontime="+86" swimtime="00:01:16.40" resultid="43968" heatid="44924" lane="2" entrytime="00:01:12.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="561" reactiontime="+84" swimtime="00:02:54.51" resultid="43969" heatid="44974" lane="5" entrytime="00:02:45.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                    <SPLIT distance="100" swimtime="00:01:21.33" />
                    <SPLIT distance="150" swimtime="00:02:12.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="663" reactiontime="+66" swimtime="00:00:35.56" resultid="43970" heatid="45027" lane="2" entrytime="00:00:36.54" entrycourse="LCM" />
                <RESULT eventid="2430" points="583" reactiontime="+78" swimtime="00:00:31.66" resultid="43971" heatid="45072" lane="7" entrytime="00:00:31.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Liliana Elisabete" lastname="Baptista" birthdate="1978-08-17" gender="F" nation="POR" license="120495" swrid="4638599" athleteid="43842">
              <RESULTS>
                <RESULT eventid="2203" points="615" reactiontime="+76" swimtime="00:01:22.40" resultid="43843" heatid="44883" lane="7" entrytime="00:01:24.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2338" points="630" reactiontime="+86" swimtime="00:00:34.22" resultid="43844" heatid="44891" lane="4" entrytime="00:00:36.15" entrycourse="LCM" />
                <RESULT eventid="2308" points="612" reactiontime="+82" swimtime="00:03:01.28" resultid="43845" heatid="44915" lane="7" entrytime="00:03:09.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                    <SPLIT distance="100" swimtime="00:01:26.90" />
                    <SPLIT distance="150" swimtime="00:02:13.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="646" reactiontime="+108" swimtime="00:00:36.63" resultid="43846" heatid="45027" lane="8" entrytime="00:00:38.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Trigueiros" lastname="Cunha" birthdate="1964-03-27" gender="F" nation="POR" license="132357" swrid="5065800" athleteid="43863">
              <RESULTS>
                <RESULT eventid="2607" points="389" reactiontime="+110" swimtime="00:00:51.76" resultid="43864" heatid="45099" lane="3" entrytime="00:00:51.83" entrycourse="LCM" />
                <RESULT eventid="2637" points="379" reactiontime="+116" swimtime="00:01:27.93" resultid="43865" heatid="44954" lane="7" entrytime="00:01:32.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="305" reactiontime="+104" swimtime="00:07:11.91" resultid="43866" heatid="45009" lane="4" entrytime="00:07:37.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.11" />
                    <SPLIT distance="100" swimtime="00:01:37.26" />
                    <SPLIT distance="150" swimtime="00:02:31.35" />
                    <SPLIT distance="200" swimtime="00:03:27.81" />
                    <SPLIT distance="250" swimtime="00:04:25.24" />
                    <SPLIT distance="300" swimtime="00:05:22.93" />
                    <SPLIT distance="350" swimtime="00:06:18.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" status="DNS" swimtime="00:00:00.00" resultid="43867" heatid="45120" lane="1" entrytime="00:01:55.56" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GDNFAMA" nation="POR" region="ANNP" clubid="42378" swrid="65898" name="Grupo Desp. Natacao V. N. Famalicao" shortname="Famalicao">
          <ATHLETES>
            <ATHLETE firstname="Antonio Sergio" lastname="Costa" birthdate="1984-03-23" gender="M" nation="POR" license="214235" swrid="4564417" athleteid="43805">
              <RESULTS>
                <RESULT eventid="2622" points="510" reactiontime="+85" swimtime="00:03:09.37" resultid="43806" heatid="44878" lane="4" entrytime="00:02:59.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                    <SPLIT distance="100" swimtime="00:01:25.88" />
                    <SPLIT distance="150" swimtime="00:02:15.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="500" reactiontime="+86" swimtime="00:00:36.79" resultid="43807" heatid="44948" lane="8" entrytime="00:00:38.20" />
                <RESULT eventid="2445" points="526" reactiontime="+89" swimtime="00:01:22.32" resultid="43808" heatid="44998" lane="4" entrytime="00:01:19.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Emanuel" lastname="Vaz" birthdate="1991-06-04" gender="M" nation="POR" license="15628" swrid="4269379" athleteid="43825">
              <RESULTS>
                <RESULT eventid="2263" points="706" reactiontime="+81" swimtime="00:04:39.09" resultid="43826" heatid="45131" lane="4" entrytime="00:04:10.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                    <SPLIT distance="100" swimtime="00:01:04.52" />
                    <SPLIT distance="150" swimtime="00:01:39.19" />
                    <SPLIT distance="200" swimtime="00:02:14.32" />
                    <SPLIT distance="250" swimtime="00:02:50.51" />
                    <SPLIT distance="300" swimtime="00:03:26.37" />
                    <SPLIT distance="350" swimtime="00:04:02.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jorge Manuel" lastname="Maia" birthdate="1989-05-02" gender="M" nation="POR" license="23220" swrid="4061673" athleteid="43817">
              <RESULTS>
                <RESULT eventid="2682" points="757" reactiontime="+72" swimtime="00:00:27.45" resultid="43818" heatid="44901" lane="3" entrytime="00:00:27.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helio Joaquim" lastname="Machado" birthdate="1983-03-09" gender="M" nation="POR" license="214217" athleteid="43815">
              <RESULTS>
                <RESULT eventid="1058" points="223" swimtime="00:14:42.47" resultid="43816" heatid="45079" lane="5" entrytime="00:18:15.27">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.36" />
                    <SPLIT distance="200" swimtime="00:03:30.82" />
                    <SPLIT distance="300" swimtime="00:05:21.76" />
                    <SPLIT distance="400" swimtime="00:07:16.75" />
                    <SPLIT distance="500" swimtime="00:09:10.05" />
                    <SPLIT distance="600" swimtime="00:11:01.32" />
                    <SPLIT distance="700" swimtime="00:12:53.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nuno Miguel" lastname="Macedo" birthdate="1982-06-29" gender="M" nation="POR" license="23308" swrid="4061678" athleteid="43811">
              <RESULTS>
                <RESULT eventid="2188" points="547" reactiontime="+72" swimtime="00:00:35.71" resultid="43812" heatid="44947" lane="4" entrytime="00:00:38.45" />
                <RESULT eventid="2415" points="510" reactiontime="+74" swimtime="00:01:05.03" resultid="43813" heatid="45113" lane="5" entrytime="00:01:03.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="551" reactiontime="+78" swimtime="00:00:28.70" resultid="43814" heatid="45045" lane="3" entrytime="00:00:27.90" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Jose" lastname="Ferreira" birthdate="1965-06-10" gender="M" nation="POR" license="214216" athleteid="43809">
              <RESULTS>
                <RESULT eventid="1058" points="176" swimtime="00:16:51.22" resultid="43810" heatid="45079" lane="3" entrytime="00:18:16.35">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.71" />
                    <SPLIT distance="200" swimtime="00:03:53.41" />
                    <SPLIT distance="300" swimtime="00:06:03.29" />
                    <SPLIT distance="400" swimtime="00:08:13.80" />
                    <SPLIT distance="500" swimtime="00:10:24.20" />
                    <SPLIT distance="600" swimtime="00:12:32.37" />
                    <SPLIT distance="700" swimtime="00:14:40.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adriano Miguel" lastname="Niz" birthdate="1986-03-05" gender="M" nation="POR" license="23013" swrid="4064351" athleteid="43819">
              <RESULTS>
                <RESULT comment="Rec Nac Esc C" eventid="2622" points="815" reactiontime="+81" swimtime="00:02:42.04" resultid="43820" heatid="44879" lane="5" entrytime="00:02:38.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="100" swimtime="00:01:17.57" />
                    <SPLIT distance="150" swimtime="00:02:00.02" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rec Nac Esc C" eventid="2218" points="1002" reactiontime="+71" swimtime="00:02:13.11" resultid="43821" heatid="44921" lane="4" entrytime="00:02:10.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:06.30" />
                    <SPLIT distance="150" swimtime="00:01:40.15" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rec Nac Esc C" eventid="2385" points="810" reactiontime="+79" swimtime="00:02:21.69" resultid="43822" heatid="44982" lane="4" entrytime="00:02:17.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.41" />
                    <SPLIT distance="100" swimtime="00:01:05.09" />
                    <SPLIT distance="150" swimtime="00:01:46.97" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rec Nac Esc C" eventid="2567" points="894" reactiontime="+80" swimtime="00:02:19.70" resultid="43823" heatid="45030" lane="4" entrytime="00:02:07.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                    <SPLIT distance="100" swimtime="00:01:04.35" />
                    <SPLIT distance="150" swimtime="00:01:40.61" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rec Nac Esc C" eventid="2248" points="769" reactiontime="+83" swimtime="00:05:11.00" resultid="43824" heatid="45062" lane="4" entrytime="00:04:30.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                    <SPLIT distance="100" swimtime="00:01:05.86" />
                    <SPLIT distance="150" swimtime="00:01:43.62" />
                    <SPLIT distance="200" swimtime="00:02:21.40" />
                    <SPLIT distance="250" swimtime="00:03:06.18" />
                    <SPLIT distance="300" swimtime="00:03:51.10" />
                    <SPLIT distance="350" swimtime="00:04:28.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="00617" nation="ESP" region="11115" clubid="41516" swrid="67768" name="A.D. Fogar">
          <ATHLETES>
            <ATHLETE firstname="Elisa" lastname="Pichel Garcia" birthdate="1984-05-16" gender="F" nation="ESP" license="1037385" swrid="5312633" athleteid="41522">
              <RESULTS>
                <RESULT eventid="2338" status="WDR" swimtime="00:00:00.00" resultid="41523" entrytime="00:00:33.69" entrycourse="SCM" />
                <RESULT eventid="2278" status="WDR" swimtime="00:00:00.00" resultid="41524" entrytime="00:02:22.87" entrycourse="SCM" />
                <RESULT eventid="2637" status="WDR" swimtime="00:00:00.00" resultid="41525" entrytime="00:01:08.86" entrycourse="SCM" />
                <RESULT eventid="2430" status="WDR" swimtime="00:00:00.00" resultid="41526" entrytime="00:00:30.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Josue" lastname="Pantoja Guio" birthdate="1978-05-02" gender="M" nation="ESP" license="1050717" swrid="5208883" athleteid="41517">
              <RESULTS>
                <RESULT eventid="2682" status="WDR" swimtime="00:00:00.00" resultid="41518" entrytime="00:00:29.76" entrycourse="SCM" />
                <RESULT eventid="2507" status="WDR" swimtime="00:00:00.00" resultid="41519" entrytime="00:02:17.83" entrycourse="SCM" />
                <RESULT eventid="2415" status="WDR" swimtime="00:00:00.00" resultid="41520" entrytime="00:00:58.88" />
                <RESULT eventid="2652" status="WDR" swimtime="00:00:00.00" resultid="41521" entrytime="00:00:28.10" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="VKGS" nation="POR" region="ANL" clubid="42992" swrid="75140" name="Vikings Sports Club" shortname="Vikings">
          <ATHLETES>
            <ATHLETE firstname="Sofia Prates" lastname="Silvestre" birthdate="1995-01-02" gender="F" nation="POR" license="121320" swrid="4691597" athleteid="42993">
              <RESULTS>
                <RESULT eventid="2552" points="662" reactiontime="+79" swimtime="00:01:11.25" resultid="42994" heatid="44924" lane="3" entrytime="00:01:08.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="668" reactiontime="+77" swimtime="00:01:05.49" resultid="42995" heatid="44957" lane="5" entrytime="00:01:01.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="723" reactiontime="+77" swimtime="00:05:00.65" resultid="42996" heatid="45013" lane="5" entrytime="00:05:06.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="100" swimtime="00:01:07.50" />
                    <SPLIT distance="150" swimtime="00:01:45.73" />
                    <SPLIT distance="200" swimtime="00:02:24.78" />
                    <SPLIT distance="250" swimtime="00:03:04.02" />
                    <SPLIT distance="300" swimtime="00:03:43.13" />
                    <SPLIT distance="350" swimtime="00:04:22.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="651" reactiontime="+75" swimtime="00:00:30.11" resultid="42997" heatid="45073" lane="5" entrytime="00:00:28.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CNV" nation="POR" region="ANNP" clubid="42919" swrid="76517" name="Clube de Natacao de Valongo" shortname="Natacao de Valongo">
          <ATHLETES>
            <ATHLETE firstname="Luis Miguel" lastname="Nunes" birthdate="1974-10-03" gender="M" nation="POR" license="209668" swrid="5344123" athleteid="43997">
              <RESULTS>
                <RESULT eventid="2293" status="DNS" swimtime="00:00:00.00" resultid="43998" heatid="45017" lane="7" entrytime="00:00:47.47" entrycourse="SCM" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="43999" heatid="45037" lane="4" entrytime="00:00:34.82" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor Manuel" lastname="Cardoso" birthdate="1972-12-02" gender="M" nation="POR" license="207728" swrid="4885761" athleteid="43987">
              <RESULTS>
                <RESULT eventid="1058" points="286" swimtime="00:13:23.82" resultid="43988" heatid="45081" lane="3" entrytime="00:14:09.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.47" />
                    <SPLIT distance="200" swimtime="00:03:12.84" />
                    <SPLIT distance="300" swimtime="00:04:57.36" />
                    <SPLIT distance="400" swimtime="00:06:42.55" />
                    <SPLIT distance="500" swimtime="00:08:25.99" />
                    <SPLIT distance="600" swimtime="00:10:08.23" />
                    <SPLIT distance="700" swimtime="00:11:50.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="284" reactiontime="+85" swimtime="00:00:40.37" resultid="43989" heatid="44894" lane="4" entrytime="00:00:40.47" entrycourse="LCM" />
                <RESULT eventid="2188" points="312" reactiontime="+86" swimtime="00:00:44.04" resultid="43990" heatid="44945" lane="6" entrytime="00:00:42.33" entrycourse="SCM" />
                <RESULT eventid="2415" points="377" reactiontime="+72" swimtime="00:01:17.29" resultid="43991" heatid="45109" lane="8" entrytime="00:01:16.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="424" reactiontime="+76" swimtime="00:00:33.08" resultid="43992" heatid="45037" lane="8" entrytime="00:00:36.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Attila Janus" lastname="Ambrus" birthdate="1974-05-16" gender="M" nation="POR" license="213595" swrid="5451866" athleteid="43983">
              <RESULTS>
                <RESULT eventid="1058" status="WDR" swimtime="00:00:00.00" resultid="43984" entrytime="00:15:10.00" />
                <RESULT eventid="2682" status="WDR" swimtime="00:00:00.00" resultid="43985" entrytime="00:00:55.00" />
                <RESULT eventid="2415" status="WDR" swimtime="00:00:00.00" resultid="43986" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo Jorge" lastname="Fernandes" birthdate="1972-06-14" gender="M" nation="POR" license="14684" swrid="4574788" athleteid="43993">
              <RESULTS>
                <RESULT eventid="2537" status="WDR" swimtime="00:00:00.00" resultid="43994" entrytime="00:01:30.25" entrycourse="SCM" />
                <RESULT eventid="2682" status="WDR" swimtime="00:00:00.00" resultid="43995" entrytime="00:00:36.47" entrycourse="LCM" />
                <RESULT eventid="2263" status="WDR" swimtime="00:00:00.00" resultid="43996" entrytime="00:06:18.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelo Porto" lastname="Rodrigues" birthdate="1982-03-15" gender="M" nation="POR" license="205613" swrid="5260608" athleteid="44006">
              <RESULTS>
                <RESULT eventid="2188" points="415" reactiontime="+76" swimtime="00:00:39.15" resultid="44007" heatid="44948" lane="7" entrytime="00:00:38.07" entrycourse="LCM" />
                <RESULT eventid="2385" points="436" reactiontime="+84" swimtime="00:02:54.18" resultid="44008" heatid="44980" lane="1" entrytime="00:02:54.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                    <SPLIT distance="100" swimtime="00:01:23.30" />
                    <SPLIT distance="150" swimtime="00:02:13.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="434" reactiontime="+89" swimtime="00:05:38.70" resultid="44009" heatid="45129" lane="8" entrytime="00:05:53.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                    <SPLIT distance="100" swimtime="00:01:17.41" />
                    <SPLIT distance="150" swimtime="00:01:59.79" />
                    <SPLIT distance="200" swimtime="00:02:43.00" />
                    <SPLIT distance="250" swimtime="00:03:26.97" />
                    <SPLIT distance="300" swimtime="00:04:11.37" />
                    <SPLIT distance="350" swimtime="00:04:56.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="464" reactiontime="+85" swimtime="00:00:30.39" resultid="44010" heatid="45039" lane="2" entrytime="00:00:33.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Susana Maria" lastname="Soares" birthdate="1970-02-19" gender="F" nation="POR" license="26158" swrid="4575644" athleteid="44011">
              <RESULTS>
                <RESULT eventid="1060" points="203" swimtime="00:16:46.85" resultid="44012" heatid="45075" lane="6" entrytime="00:16:45.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.38" />
                    <SPLIT distance="200" swimtime="00:03:59.84" />
                    <SPLIT distance="300" swimtime="00:06:07.84" />
                    <SPLIT distance="400" swimtime="00:08:16.81" />
                    <SPLIT distance="500" swimtime="00:10:25.91" />
                    <SPLIT distance="600" swimtime="00:12:34.09" />
                    <SPLIT distance="700" swimtime="00:14:43.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="363" reactiontime="+97" swimtime="00:00:51.45" resultid="44013" heatid="45100" lane="1" entrytime="00:00:50.00" />
                <RESULT eventid="2637" points="232" reactiontime="+109" swimtime="00:01:42.85" resultid="44014" heatid="44953" lane="1" entrytime="00:01:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="379" reactiontime="+100" swimtime="00:01:54.62" resultid="44015" heatid="45119" lane="3" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="226" reactiontime="+105" swimtime="00:07:52.84" resultid="44016" heatid="45009" lane="8" entrytime="00:08:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.61" />
                    <SPLIT distance="100" swimtime="00:01:47.16" />
                    <SPLIT distance="150" swimtime="00:02:47.66" />
                    <SPLIT distance="200" swimtime="00:03:48.88" />
                    <SPLIT distance="250" swimtime="00:04:51.52" />
                    <SPLIT distance="300" swimtime="00:05:54.77" />
                    <SPLIT distance="350" swimtime="00:06:55.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago Melo" lastname="Pereira" birthdate="1979-01-29" gender="M" nation="POR" license="208402" swrid="5326901" athleteid="44000">
              <RESULTS>
                <RESULT eventid="2682" status="DNS" swimtime="00:00:00.00" resultid="44001" heatid="44893" lane="3" entrytime="00:00:50.00" />
                <RESULT eventid="2188" points="447" reactiontime="+80" swimtime="00:00:39.88" resultid="44002" heatid="44943" lane="2" entrytime="00:00:45.00" />
                <RESULT comment="403 - Falsa partida - SW 4.4" eventid="2385" reactiontime="+84" status="DSQ" swimtime="00:03:26.47" resultid="44003" heatid="44978" lane="8" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                    <SPLIT distance="100" swimtime="00:01:41.57" />
                    <SPLIT distance="150" swimtime="00:02:36.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="235" reactiontime="+82" swimtime="00:00:45.99" resultid="44004" heatid="45016" lane="6" entrytime="00:00:51.23" entrycourse="SCM" />
                <RESULT eventid="2652" points="295" reactiontime="+93" swimtime="00:00:36.89" resultid="44005" heatid="45037" lane="1" entrytime="00:00:36.15" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CNF" nation="POR" region="ANMAD" clubid="43172" swrid="65893" name="Clube Naval do Funchal" shortname="Naval do Funchal">
          <ATHLETES>
            <ATHLETE firstname="Joao Pedro" lastname="Sousa" birthdate="1974-06-29" gender="M" nation="POR" license="128627" swrid="4931932" athleteid="43173">
              <RESULTS>
                <RESULT eventid="2507" points="649" reactiontime="+73" swimtime="00:02:17.85" resultid="43174" heatid="45096" lane="7" entrytime="00:02:15.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.23" />
                    <SPLIT distance="100" swimtime="00:01:06.63" />
                    <SPLIT distance="150" swimtime="00:01:42.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="763" reactiontime="+79" swimtime="00:01:01.10" resultid="43175" heatid="45114" lane="6" entrytime="00:01:02.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="620" reactiontime="+76" swimtime="00:05:00.38" resultid="43176" heatid="45131" lane="2" entrytime="00:04:54.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:09.19" />
                    <SPLIT distance="150" swimtime="00:01:46.91" />
                    <SPLIT distance="200" swimtime="00:02:25.63" />
                    <SPLIT distance="250" swimtime="00:03:04.30" />
                    <SPLIT distance="300" swimtime="00:03:43.62" />
                    <SPLIT distance="350" swimtime="00:04:22.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="697" reactiontime="+68" swimtime="00:00:28.04" resultid="43177" heatid="45044" lane="5" entrytime="00:00:28.63" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCP" nation="POR" region="ANL" clubid="41931" swrid="72842" name="Sporting Clube de Portugal" shortname="Sporting">
          <ATHLETES>
            <ATHLETE firstname="Helena Paula" lastname="Carvalho" birthdate="1964-05-03" gender="F" nation="POR" license="17549" swrid="4800234" athleteid="42966">
              <RESULTS>
                <RESULT eventid="2173" points="599" swimtime="00:03:44.58" resultid="42967" heatid="45089" lane="8" entrytime="00:03:41.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.08" />
                    <SPLIT distance="100" swimtime="00:01:48.94" />
                    <SPLIT distance="150" swimtime="00:02:47.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="430" reactiontime="+107" swimtime="00:00:50.05" resultid="42968" heatid="45100" lane="5" entrytime="00:00:48.98" entrycourse="LCM" />
                <RESULT eventid="2460" points="494" reactiontime="+102" swimtime="00:01:47.23" resultid="42969" heatid="45121" lane="8" entrytime="00:01:48.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="338" reactiontime="+101" swimtime="00:06:57.09" resultid="42970" heatid="45011" lane="4" entrytime="00:06:29.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.17" />
                    <SPLIT distance="100" swimtime="00:01:39.57" />
                    <SPLIT distance="150" swimtime="00:02:32.45" />
                    <SPLIT distance="200" swimtime="00:03:26.25" />
                    <SPLIT distance="250" swimtime="00:04:20.20" />
                    <SPLIT distance="300" swimtime="00:05:13.54" />
                    <SPLIT distance="350" swimtime="00:06:06.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Miguel" lastname="Batalha" birthdate="1976-12-18" gender="M" nation="POR" license="202103" swrid="5197027" athleteid="42960">
              <RESULTS>
                <RESULT eventid="2682" points="557" reactiontime="+87" swimtime="00:00:32.27" resultid="42961" heatid="44898" lane="6" entrytime="00:00:31.43" entrycourse="LCM" />
                <RESULT eventid="2188" points="449" reactiontime="+84" swimtime="00:00:39.02" resultid="42962" heatid="44948" lane="1" entrytime="00:00:38.08" entrycourse="LCM" />
                <RESULT eventid="2415" points="520" reactiontime="+87" swimtime="00:01:09.43" resultid="42963" heatid="45113" lane="1" entrytime="00:01:04.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="429" reactiontime="+88" swimtime="00:01:31.30" resultid="42964" heatid="44996" lane="6" entrytime="00:01:32.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="573" reactiontime="+91" swimtime="00:00:29.94" resultid="42965" heatid="45043" lane="1" entrytime="00:00:29.29" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo Paula" lastname="Carvalho" birthdate="1961-03-23" gender="M" nation="POR" license="25645" swrid="4574562" athleteid="42971">
              <RESULTS>
                <RESULT comment="Rec Nac Esc H" eventid="1058" points="916" swimtime="00:10:44.28" resultid="42972" heatid="45085" lane="2" entrytime="00:10:50.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.54" />
                    <SPLIT distance="200" swimtime="00:02:38.31" />
                    <SPLIT distance="300" swimtime="00:04:00.18" />
                    <SPLIT distance="400" swimtime="00:05:20.99" />
                    <SPLIT distance="500" swimtime="00:06:42.61" />
                    <SPLIT distance="600" swimtime="00:08:03.98" />
                    <SPLIT distance="700" swimtime="00:09:25.08" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rec Nac Esc H" eventid="2218" points="925" reactiontime="+72" swimtime="00:02:47.34" resultid="42973" heatid="44921" lane="6" entrytime="00:02:31.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.31" />
                    <SPLIT distance="100" swimtime="00:01:22.01" />
                    <SPLIT distance="150" swimtime="00:02:05.48" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rec Nac Esc H" eventid="2385" points="896" reactiontime="+89" swimtime="00:02:44.91" resultid="42974" heatid="44982" lane="2" entrytime="00:02:34.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                    <SPLIT distance="100" swimtime="00:01:15.58" />
                    <SPLIT distance="150" swimtime="00:02:07.11" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rec Nac Esc H" eventid="2567" points="1132" reactiontime="+89" swimtime="00:02:42.35" resultid="42975" heatid="45030" lane="3" entrytime="00:02:36.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:15.53" />
                    <SPLIT distance="150" swimtime="00:01:57.24" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rec Nac Esc H" eventid="2248" points="900" reactiontime="+85" swimtime="00:05:58.46" resultid="42976" heatid="45062" lane="7" entrytime="00:05:41.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                    <SPLIT distance="100" swimtime="00:01:11.52" />
                    <SPLIT distance="150" swimtime="00:02:01.79" />
                    <SPLIT distance="200" swimtime="00:02:49.83" />
                    <SPLIT distance="250" swimtime="00:03:45.03" />
                    <SPLIT distance="300" swimtime="00:04:40.23" />
                    <SPLIT distance="350" swimtime="00:05:20.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Samuel" lastname="Duarte" birthdate="1965-03-11" gender="M" nation="POR" license="120465" swrid="4638597" athleteid="42977">
              <RESULTS>
                <RESULT eventid="2622" status="DNS" swimtime="00:00:00.00" resultid="42978" heatid="44879" lane="2" entrytime="00:02:48.40" entrycourse="LCM" />
                <RESULT eventid="2188" status="DNS" swimtime="00:00:00.00" resultid="42979" heatid="44950" lane="7" entrytime="00:00:34.26" entrycourse="LCM" />
                <RESULT eventid="2445" status="DNS" swimtime="00:00:00.00" resultid="42980" heatid="44999" lane="6" entrytime="00:01:15.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hugo Andre" lastname="Afonso" birthdate="1976-12-23" gender="M" nation="POR" license="204884" swrid="5216335" athleteid="42954">
              <RESULTS>
                <RESULT eventid="1058" points="390" swimtime="00:12:05.45" resultid="42955" heatid="45083" lane="2" entrytime="00:12:43.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.85" />
                    <SPLIT distance="200" swimtime="00:02:57.15" />
                    <SPLIT distance="300" swimtime="00:04:29.56" />
                    <SPLIT distance="400" swimtime="00:06:02.59" />
                    <SPLIT distance="500" swimtime="00:07:35.15" />
                    <SPLIT distance="600" swimtime="00:09:06.53" />
                    <SPLIT distance="700" swimtime="00:10:37.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="428" reactiontime="+90" swimtime="00:01:14.11" resultid="42956" heatid="45109" lane="3" entrytime="00:01:14.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="394" reactiontime="+91" swimtime="00:05:49.41" resultid="42957" heatid="45129" lane="3" entrytime="00:05:45.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                    <SPLIT distance="100" swimtime="00:01:20.00" />
                    <SPLIT distance="150" swimtime="00:02:04.99" />
                    <SPLIT distance="200" swimtime="00:02:50.78" />
                    <SPLIT distance="250" swimtime="00:03:36.93" />
                    <SPLIT distance="300" swimtime="00:04:22.15" />
                    <SPLIT distance="350" swimtime="00:05:07.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="449" reactiontime="+87" swimtime="00:00:32.46" resultid="42958" heatid="45038" lane="4" entrytime="00:00:33.89" entrycourse="LCM" />
                <RESULT eventid="2507" points="363" reactiontime="+87" swimtime="00:02:47.25" resultid="42959" heatid="45092" lane="4" entrytime="00:02:52.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                    <SPLIT distance="100" swimtime="00:01:18.60" />
                    <SPLIT distance="150" swimtime="00:02:03.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patrick" lastname="Santos" birthdate="1979-07-22" gender="M" nation="POR" license="26609" swrid="4575768" athleteid="42986">
              <RESULTS>
                <RESULT eventid="1058" points="562" swimtime="00:10:37.66" resultid="42987" heatid="45085" lane="6" entrytime="00:10:30.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.92" />
                    <SPLIT distance="200" swimtime="00:02:37.21" />
                    <SPLIT distance="300" swimtime="00:03:57.04" />
                    <SPLIT distance="400" swimtime="00:05:17.59" />
                    <SPLIT distance="500" swimtime="00:06:38.29" />
                    <SPLIT distance="600" swimtime="00:07:58.95" />
                    <SPLIT distance="700" swimtime="00:09:18.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2622" points="605" reactiontime="+83" swimtime="00:02:58.32" resultid="42988" heatid="44879" lane="1" entrytime="00:02:51.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                    <SPLIT distance="100" swimtime="00:01:25.36" />
                    <SPLIT distance="150" swimtime="00:02:12.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="528" reactiontime="+81" swimtime="00:02:43.75" resultid="42989" heatid="44981" lane="4" entrytime="00:02:38.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                    <SPLIT distance="100" swimtime="00:01:20.69" />
                    <SPLIT distance="150" swimtime="00:02:05.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" points="469" reactiontime="+82" swimtime="00:02:50.27" resultid="42990" heatid="45030" lane="6" entrytime="00:02:38.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                    <SPLIT distance="100" swimtime="00:01:20.33" />
                    <SPLIT distance="150" swimtime="00:02:04.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="555" reactiontime="+83" swimtime="00:05:44.26" resultid="42991" heatid="45062" lane="6" entrytime="00:05:31.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                    <SPLIT distance="100" swimtime="00:01:17.64" />
                    <SPLIT distance="150" swimtime="00:02:06.41" />
                    <SPLIT distance="200" swimtime="00:02:53.09" />
                    <SPLIT distance="250" swimtime="00:03:39.55" />
                    <SPLIT distance="300" swimtime="00:04:26.27" />
                    <SPLIT distance="350" swimtime="00:05:05.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jorge Sequeira" lastname="Lima" birthdate="1967-07-27" gender="M" nation="POR" license="10524" swrid="5125094" athleteid="42981">
              <RESULTS>
                <RESULT eventid="2622" points="594" reactiontime="+91" swimtime="00:03:10.37" resultid="42982" heatid="44878" lane="3" entrytime="00:03:05.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.84" />
                    <SPLIT distance="100" swimtime="00:01:30.85" />
                    <SPLIT distance="150" swimtime="00:02:22.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="397" reactiontime="+98" swimtime="00:02:53.11" resultid="42983" heatid="45094" lane="1" entrytime="00:02:39.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.13" />
                    <SPLIT distance="100" swimtime="00:01:24.13" />
                    <SPLIT distance="150" swimtime="00:02:10.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="517" reactiontime="+79" swimtime="00:00:38.77" resultid="42984" heatid="44948" lane="6" entrytime="00:00:37.85" entrycourse="LCM" />
                <RESULT eventid="2445" points="562" reactiontime="+88" swimtime="00:01:27.80" resultid="42985" heatid="44997" lane="3" entrytime="00:01:27.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GCVR" nation="POR" region="ARNN" clubid="42999" swrid="66442" name="Ginasio Clube de Vila Real" shortname="Ginasio de Vila Real">
          <ATHLETES>
            <ATHLETE firstname="Daniel Pinto" lastname="Conceicao" birthdate="1994-10-06" gender="M" nation="POR" license="123283" swrid="4756547" athleteid="43000">
              <RESULTS>
                <RESULT eventid="2682" status="DNS" swimtime="00:00:00.00" resultid="43001" heatid="44897" lane="8" entrytime="00:00:35.18" entrycourse="LCM" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="43002" heatid="45043" lane="8" entrytime="00:00:29.47" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alessia Santos" lastname="Teixeira" birthdate="1995-06-21" gender="F" nation="POR" license="207255" swrid="5287899" athleteid="43007">
              <RESULTS>
                <RESULT eventid="2338" points="380" reactiontime="+81" swimtime="00:00:38.37" resultid="43008" heatid="44891" lane="7" entrytime="00:00:37.87" entrycourse="LCM" />
                <RESULT eventid="2460" points="413" reactiontime="+72" swimtime="00:01:37.11" resultid="43009" heatid="45123" lane="2" entrytime="00:01:30.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="417" reactiontime="+75" swimtime="00:00:34.91" resultid="43010" heatid="45070" lane="1" entrytime="00:00:36.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raul Morais" lastname="Santos" birthdate="1969-10-14" gender="M" nation="POR" license="127870" swrid="4905850" athleteid="43005">
              <RESULTS>
                <RESULT eventid="2652" points="458" reactiontime="+77" swimtime="00:00:32.58" resultid="43006" heatid="45041" lane="1" entrytime="00:00:31.26" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Pereira" lastname="Matos" birthdate="1983-06-23" gender="M" nation="POR" license="24788" swrid="4073985" athleteid="43003">
              <RESULTS>
                <RESULT eventid="2652" points="601" reactiontime="+84" swimtime="00:00:27.87" resultid="43004" heatid="45047" lane="4" entrytime="00:00:26.45" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="UDO" nation="POR" region="ANCNP" clubid="41774" swrid="71292" name="Uniao Desportiva Oliveirense" shortname="UD Oliveirense">
          <ATHLETES>
            <ATHLETE firstname="Jose Pedro" lastname="Bernardes" birthdate="1995-06-30" gender="M" nation="POR" license="110572" swrid="4375288" athleteid="43600">
              <RESULTS>
                <RESULT eventid="2263" points="440" reactiontime="+98" swimtime="00:05:29.68" resultid="43601" heatid="45130" lane="7" entrytime="00:05:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:01:18.22" />
                    <SPLIT distance="150" swimtime="00:02:00.96" />
                    <SPLIT distance="200" swimtime="00:02:43.39" />
                    <SPLIT distance="250" swimtime="00:03:25.31" />
                    <SPLIT distance="300" swimtime="00:04:06.81" />
                    <SPLIT distance="350" swimtime="00:04:49.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="487" reactiontime="+73" swimtime="00:00:34.03" resultid="43602" heatid="45022" lane="2" entrytime="00:00:31.50" />
                <RESULT eventid="2248" status="DNS" swimtime="00:00:00.00" resultid="43603" heatid="45061" lane="2" entrytime="00:06:25.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco Nunes" lastname="Silva" birthdate="1995-03-18" gender="M" nation="POR" license="123546" swrid="4756723" athleteid="43604">
              <RESULTS>
                <RESULT eventid="2293" points="415" reactiontime="+67" swimtime="00:00:35.88" resultid="43605" heatid="45020" lane="4" entrytime="00:00:33.50" />
                <RESULT eventid="2652" points="519" reactiontime="+72" swimtime="00:00:28.80" resultid="43606" heatid="45045" lane="6" entrytime="00:00:28.00" />
                <RESULT eventid="2248" points="374" reactiontime="+75" swimtime="00:06:36.06" resultid="43607" heatid="45060" lane="5" entrytime="00:06:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                    <SPLIT distance="100" swimtime="00:01:22.32" />
                    <SPLIT distance="150" swimtime="00:02:16.75" />
                    <SPLIT distance="200" swimtime="00:03:09.90" />
                    <SPLIT distance="250" swimtime="00:04:07.15" />
                    <SPLIT distance="300" swimtime="00:05:05.47" />
                    <SPLIT distance="350" swimtime="00:05:52.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aleksandro" lastname="Aita" birthdate="1974-06-13" gender="M" nation="BRA" license="214136" swrid="5467363" athleteid="43596">
              <RESULTS>
                <RESULT eventid="1058" points="424" swimtime="00:11:45.56" resultid="43597" heatid="45084" lane="2" entrytime="00:11:40.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.84" />
                    <SPLIT distance="200" swimtime="00:02:46.75" />
                    <SPLIT distance="300" swimtime="00:04:14.77" />
                    <SPLIT distance="400" swimtime="00:05:44.51" />
                    <SPLIT distance="500" swimtime="00:07:14.89" />
                    <SPLIT distance="600" swimtime="00:08:46.29" />
                    <SPLIT distance="700" swimtime="00:10:17.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="418" reactiontime="+76" swimtime="00:00:39.98" resultid="43598" heatid="44949" lane="7" entrytime="00:00:36.00" />
                <RESULT eventid="2263" points="409" reactiontime="+88" swimtime="00:05:45.14" resultid="43599" heatid="45127" lane="5" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                    <SPLIT distance="100" swimtime="00:01:21.16" />
                    <SPLIT distance="150" swimtime="00:02:04.94" />
                    <SPLIT distance="200" swimtime="00:02:48.99" />
                    <SPLIT distance="250" swimtime="00:03:33.70" />
                    <SPLIT distance="300" swimtime="00:04:18.20" />
                    <SPLIT distance="350" swimtime="00:05:02.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CFP" nation="POR" region="ANNP" clubid="41927" swrid="65888" name="Clube Fluvial Portuense" shortname="Fluvial Portuense">
          <ATHLETES>
            <ATHLETE firstname="Luis Manuel" lastname="Sousa" birthdate="1966-12-10" gender="M" nation="POR" license="14630" swrid="4575928" athleteid="43550">
              <RESULTS>
                <RESULT eventid="2263" points="377" reactiontime="+93" swimtime="00:06:22.41" resultid="43551" heatid="45127" lane="6" entrytime="00:06:35.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                    <SPLIT distance="100" swimtime="00:01:25.09" />
                    <SPLIT distance="150" swimtime="00:02:14.73" />
                    <SPLIT distance="200" swimtime="00:03:04.43" />
                    <SPLIT distance="250" swimtime="00:03:55.37" />
                    <SPLIT distance="300" swimtime="00:04:45.06" />
                    <SPLIT distance="350" swimtime="00:05:35.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="325" reactiontime="+75" swimtime="00:00:45.51" resultid="43552" heatid="45017" lane="2" entrytime="00:00:46.89" entrycourse="LCM" />
                <RESULT eventid="2652" points="517" reactiontime="+78" swimtime="00:00:33.14" resultid="43553" heatid="45038" lane="2" entrytime="00:00:34.19" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela Maria" lastname="Palhares" birthdate="1971-11-04" gender="F" nation="POR" license="209005" swrid="5322823" athleteid="43428">
              <RESULTS>
                <RESULT eventid="2203" points="396" reactiontime="+78" swimtime="00:01:42.64" resultid="43429" heatid="44882" lane="2" entrytime="00:01:37.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2278" points="346" reactiontime="+104" swimtime="00:03:16.56" resultid="43430" heatid="44902" lane="4" entrytime="00:03:31.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                    <SPLIT distance="100" swimtime="00:01:28.99" />
                    <SPLIT distance="150" swimtime="00:02:22.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="364" reactiontime="+77" swimtime="00:00:48.09" resultid="43431" heatid="45024" lane="4" entrytime="00:00:47.16" entrycourse="SCM" />
                <RESULT eventid="1060" points="340" swimtime="00:14:08.42" resultid="43432" heatid="45077" lane="7" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.54" />
                    <SPLIT distance="200" swimtime="00:03:22.89" />
                    <SPLIT distance="300" swimtime="00:05:10.81" />
                    <SPLIT distance="400" swimtime="00:07:00.76" />
                    <SPLIT distance="500" swimtime="00:08:50.04" />
                    <SPLIT distance="600" swimtime="00:10:37.74" />
                    <SPLIT distance="700" swimtime="00:12:24.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="353" reactiontime="+103" swimtime="00:06:47.92" resultid="43433" heatid="45012" lane="8" entrytime="00:06:28.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.22" />
                    <SPLIT distance="100" swimtime="00:01:34.43" />
                    <SPLIT distance="150" swimtime="00:02:27.19" />
                    <SPLIT distance="200" swimtime="00:03:19.93" />
                    <SPLIT distance="250" swimtime="00:04:12.44" />
                    <SPLIT distance="300" swimtime="00:05:05.31" />
                    <SPLIT distance="350" swimtime="00:05:58.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Paula" lastname="Dupont" birthdate="1958-07-27" gender="F" nation="POR" license="205209" swrid="5231521" athleteid="43287">
              <RESULTS>
                <RESULT eventid="1060" points="234" swimtime="00:19:07.34" resultid="43288" heatid="45074" lane="7" entrytime="00:19:28.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:06.16" />
                    <SPLIT distance="200" swimtime="00:04:25.71" />
                    <SPLIT distance="300" swimtime="00:06:52.29" />
                    <SPLIT distance="400" swimtime="00:09:19.32" />
                    <SPLIT distance="500" swimtime="00:11:45.12" />
                    <SPLIT distance="600" swimtime="00:14:12.71" />
                    <SPLIT distance="700" swimtime="00:16:41.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2173" points="369" swimtime="00:04:32.68" resultid="43289" heatid="45087" lane="1" entrytime="00:04:32.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.49" />
                    <SPLIT distance="100" swimtime="00:02:13.74" />
                    <SPLIT distance="150" swimtime="00:03:24.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="282" reactiontime="+123" swimtime="00:00:57.59" resultid="43290" heatid="45098" lane="3" entrytime="00:00:58.34" entrycourse="LCM" />
                <RESULT eventid="2460" points="301" swimtime="00:02:08.02" resultid="43291" heatid="45119" lane="8" entrytime="00:02:05.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="238" swimtime="00:09:22.79" resultid="43292" heatid="45008" lane="2" entrytime="00:09:38.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.91" />
                    <SPLIT distance="100" swimtime="00:02:11.02" />
                    <SPLIT distance="150" swimtime="00:03:22.42" />
                    <SPLIT distance="200" swimtime="00:04:34.78" />
                    <SPLIT distance="250" swimtime="00:05:48.30" />
                    <SPLIT distance="300" swimtime="00:07:00.42" />
                    <SPLIT distance="350" swimtime="00:08:12.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Ana" lastname="Fonseca" birthdate="1982-01-28" gender="F" nation="POR" license="129912" swrid="4982758" athleteid="43311">
              <RESULTS>
                <RESULT eventid="2492" points="233" reactiontime="+96" swimtime="00:07:36.39" resultid="43312" heatid="45012" lane="2" entrytime="00:06:22.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                    <SPLIT distance="100" swimtime="00:01:37.37" />
                    <SPLIT distance="150" swimtime="00:02:30.77" />
                    <SPLIT distance="200" swimtime="00:03:29.49" />
                    <SPLIT distance="250" swimtime="00:04:28.28" />
                    <SPLIT distance="300" swimtime="00:05:30.72" />
                    <SPLIT distance="350" swimtime="00:06:32.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rita Cabral" lastname="Guimaraes" birthdate="1964-12-15" gender="F" nation="POR" license="104341" swrid="5119297" athleteid="43326">
              <RESULTS>
                <RESULT eventid="1060" points="363" swimtime="00:14:07.98" resultid="43327" heatid="45077" lane="6" entrytime="00:13:24.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.31" />
                    <SPLIT distance="200" swimtime="00:03:26.52" />
                    <SPLIT distance="300" swimtime="00:05:14.87" />
                    <SPLIT distance="400" swimtime="00:07:02.31" />
                    <SPLIT distance="500" swimtime="00:08:50.48" />
                    <SPLIT distance="600" swimtime="00:10:38.11" />
                    <SPLIT distance="700" swimtime="00:12:25.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2203" points="453" reactiontime="+103" swimtime="00:01:41.73" resultid="43328" heatid="44882" lane="1" entrytime="00:01:38.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2278" points="371" swimtime="00:03:14.44" resultid="43329" heatid="44904" lane="7" entrytime="00:03:04.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.75" />
                    <SPLIT distance="100" swimtime="00:01:32.18" />
                    <SPLIT distance="150" swimtime="00:02:24.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2308" points="433" reactiontime="+85" swimtime="00:03:40.63" resultid="43330" heatid="44914" lane="6" entrytime="00:03:39.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.56" />
                    <SPLIT distance="100" swimtime="00:01:48.49" />
                    <SPLIT distance="150" swimtime="00:02:46.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="431" reactiontime="+81" swimtime="00:01:24.29" resultid="43331" heatid="44955" lane="4" entrytime="00:01:19.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Susana Maria" lastname="Lourenco" birthdate="1974-07-24" gender="F" nation="POR" license="209008" swrid="5317801" athleteid="43353">
              <RESULTS>
                <RESULT eventid="2492" points="115" swimtime="00:09:44.10" resultid="43354" heatid="45008" lane="6" entrytime="00:09:33.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.60" />
                    <SPLIT distance="100" swimtime="00:02:17.42" />
                    <SPLIT distance="150" swimtime="00:03:31.31" />
                    <SPLIT distance="200" swimtime="00:04:45.56" />
                    <SPLIT distance="250" swimtime="00:06:00.32" />
                    <SPLIT distance="300" swimtime="00:07:14.86" />
                    <SPLIT distance="350" swimtime="00:08:31.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2667" points="120" swimtime="00:05:15.24" resultid="43355" heatid="45031" lane="8" entrytime="00:04:48.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.61" />
                    <SPLIT distance="100" swimtime="00:02:29.95" />
                    <SPLIT distance="150" swimtime="00:03:52.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Luisa" lastname="Costa" birthdate="1974-05-03" gender="F" nation="POR" license="119218" swrid="4598693" athleteid="43275">
              <RESULTS>
                <RESULT eventid="1060" points="551" swimtime="00:11:47.99" resultid="43276" heatid="45078" lane="4" entrytime="00:11:11.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.12" />
                    <SPLIT distance="200" swimtime="00:02:48.86" />
                    <SPLIT distance="300" swimtime="00:04:16.55" />
                    <SPLIT distance="400" swimtime="00:05:46.30" />
                    <SPLIT distance="500" swimtime="00:07:15.64" />
                    <SPLIT distance="600" swimtime="00:08:47.09" />
                    <SPLIT distance="700" swimtime="00:10:18.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2338" points="655" reactiontime="+89" swimtime="00:00:34.74" resultid="43277" heatid="44892" lane="7" entrytime="00:00:34.26" entrycourse="LCM" />
                <RESULT eventid="2278" points="589" reactiontime="+93" swimtime="00:02:38.99" resultid="43278" heatid="44905" lane="2" entrytime="00:02:33.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                    <SPLIT distance="100" swimtime="00:01:16.36" />
                    <SPLIT distance="150" swimtime="00:01:57.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="641" reactiontime="+90" swimtime="00:02:56.30" resultid="43279" heatid="44974" lane="3" entrytime="00:02:52.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:24.26" />
                    <SPLIT distance="150" swimtime="00:02:16.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2400" points="703" reactiontime="+93" swimtime="00:06:14.04" resultid="43280" heatid="45064" lane="4" entrytime="00:05:54.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:17.06" />
                    <SPLIT distance="150" swimtime="00:02:07.87" />
                    <SPLIT distance="200" swimtime="00:02:58.36" />
                    <SPLIT distance="250" swimtime="00:03:53.22" />
                    <SPLIT distance="300" swimtime="00:04:49.09" />
                    <SPLIT distance="350" swimtime="00:05:31.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Miguel" lastname="Bernardo" birthdate="1961-04-22" gender="M" nation="POR" license="201380" swrid="5171462" athleteid="43212">
              <RESULTS>
                <RESULT eventid="2622" points="632" reactiontime="+99" swimtime="00:03:18.92" resultid="43213" heatid="44877" lane="4" entrytime="00:03:17.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.57" />
                    <SPLIT distance="100" swimtime="00:01:35.09" />
                    <SPLIT distance="150" swimtime="00:02:27.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="499" reactiontime="+94" swimtime="00:00:36.70" resultid="43214" heatid="44895" lane="5" entrytime="00:00:38.01" entrycourse="LCM" />
                <RESULT eventid="2188" points="696" reactiontime="+90" swimtime="00:00:37.99" resultid="43215" heatid="44948" lane="4" entrytime="00:00:36.97" entrycourse="LCM" />
                <RESULT eventid="2445" points="708" reactiontime="+96" swimtime="00:01:26.39" resultid="43216" heatid="44997" lane="6" entrytime="00:01:28.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="604" reactiontime="+102" swimtime="00:05:54.60" resultid="43217" heatid="45128" lane="7" entrytime="00:06:21.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.99" />
                    <SPLIT distance="100" swimtime="00:01:23.34" />
                    <SPLIT distance="150" swimtime="00:02:08.69" />
                    <SPLIT distance="200" swimtime="00:02:54.29" />
                    <SPLIT distance="250" swimtime="00:03:41.07" />
                    <SPLIT distance="300" swimtime="00:04:26.53" />
                    <SPLIT distance="350" swimtime="00:05:11.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arnaldo Silva" lastname="Martins" birthdate="1961-05-27" gender="M" nation="POR" license="129911" swrid="4982790" athleteid="43368">
              <RESULTS>
                <RESULT eventid="2445" status="DNS" swimtime="00:00:00.00" resultid="43369" heatid="44991" lane="5" entrytime="00:02:05.46" entrycourse="LCM" />
                <RESULT eventid="2385" status="DNS" swimtime="00:00:00.00" resultid="43370" heatid="44975" lane="2" entrytime="00:04:42.71" entrycourse="LCM" />
                <RESULT eventid="2263" status="DNS" swimtime="00:00:00.00" resultid="43371" heatid="45125" lane="3" entrytime="00:07:52.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Cesar" lastname="Alves" birthdate="1963-09-21" gender="M" nation="POR" license="214253" swrid="5472927" athleteid="43181">
              <RESULTS>
                <RESULT eventid="1058" points="107" swimtime="00:19:53.11" resultid="43182" heatid="45079" lane="4" entrytime="00:18:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:13.53" />
                    <SPLIT distance="200" swimtime="00:04:40.30" />
                    <SPLIT distance="300" swimtime="00:07:08.74" />
                    <SPLIT distance="400" swimtime="00:09:40.03" />
                    <SPLIT distance="500" swimtime="00:12:12.36" />
                    <SPLIT distance="600" swimtime="00:14:47.09" />
                    <SPLIT distance="700" swimtime="00:17:23.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Jorge" lastname="Marques" birthdate="1951-10-10" gender="M" nation="POR" license="130679" swrid="5001724" athleteid="43356">
              <RESULTS>
                <RESULT eventid="2622" points="277" reactiontime="+118" swimtime="00:04:55.39" resultid="43357" heatid="44873" lane="2" entrytime="00:04:44.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.76" />
                    <SPLIT distance="100" swimtime="00:02:20.77" />
                    <SPLIT distance="150" swimtime="00:03:39.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="162" reactiontime="+93" swimtime="00:00:57.84" resultid="43358" heatid="44893" lane="2" entrytime="00:00:54.68" entrycourse="LCM" />
                <RESULT eventid="2188" points="245" reactiontime="+97" swimtime="00:00:58.85" resultid="43359" heatid="44939" lane="3" entrytime="00:00:52.93" entrycourse="LCM" />
                <RESULT eventid="2293" points="211" reactiontime="+92" swimtime="00:00:58.58" resultid="43360" heatid="45014" lane="4" entrytime="00:01:02.76" entrycourse="LCM" />
                <RESULT eventid="2652" points="234" reactiontime="+91" swimtime="00:00:46.13" resultid="43361" heatid="45033" lane="5" entrytime="00:00:49.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elza Maria" lastname="Carvalho" birthdate="1976-01-13" gender="F" nation="POR" license="153144" swrid="5112926" athleteid="43238">
              <RESULTS>
                <RESULT eventid="2173" points="468" swimtime="00:03:40.08" resultid="43239" heatid="45089" lane="1" entrytime="00:03:35.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.50" />
                    <SPLIT distance="100" swimtime="00:01:44.10" />
                    <SPLIT distance="150" swimtime="00:02:41.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="491" reactiontime="+85" swimtime="00:00:45.89" resultid="43240" heatid="45101" lane="5" entrytime="00:00:44.65" entrycourse="LCM" />
                <RESULT eventid="2233" points="417" reactiontime="+104" swimtime="00:03:23.39" resultid="43241" heatid="44973" lane="8" entrytime="00:03:15.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.52" />
                    <SPLIT distance="100" swimtime="00:01:42.38" />
                    <SPLIT distance="150" swimtime="00:02:36.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="535" reactiontime="+93" swimtime="00:01:38.67" resultid="43242" heatid="45122" lane="8" entrytime="00:01:40.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2400" points="390" reactiontime="+106" swimtime="00:07:35.14" resultid="43243" heatid="45064" lane="3" entrytime="00:06:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.60" />
                    <SPLIT distance="100" swimtime="00:01:49.23" />
                    <SPLIT distance="150" swimtime="00:02:53.22" />
                    <SPLIT distance="200" swimtime="00:03:55.72" />
                    <SPLIT distance="250" swimtime="00:04:54.04" />
                    <SPLIT distance="300" swimtime="00:05:53.38" />
                    <SPLIT distance="350" swimtime="00:06:47.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Jorge" lastname="Marques" birthdate="1978-08-06" gender="M" nation="POR" license="129104" swrid="4951654" athleteid="43362">
              <RESULTS>
                <RESULT eventid="2682" points="616" reactiontime="+76" swimtime="00:00:30.43" resultid="43363" heatid="44899" lane="6" entrytime="00:00:30.33" entrycourse="LCM" />
                <RESULT eventid="2323" points="436" reactiontime="+79" swimtime="00:01:17.37" resultid="43364" heatid="44926" lane="4" entrytime="00:01:25.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="456" reactiontime="+80" swimtime="00:02:51.95" resultid="43365" heatid="44981" lane="6" entrytime="00:02:42.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:18.63" />
                    <SPLIT distance="150" swimtime="00:02:11.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="454" reactiontime="+76" swimtime="00:00:36.95" resultid="43366" heatid="45020" lane="7" entrytime="00:00:35.06" entrycourse="LCM" />
                <RESULT eventid="2652" points="631" reactiontime="+76" swimtime="00:00:28.65" resultid="43367" heatid="45046" lane="8" entrytime="00:00:27.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marilia Laura" lastname="Silva" birthdate="1952-05-01" gender="F" nation="POR" license="131783" swrid="5036833" athleteid="43533">
              <RESULTS>
                <RESULT eventid="2278" points="134" swimtime="00:05:16.69" resultid="43534" heatid="44902" lane="1" entrytime="00:05:15.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.62" />
                    <SPLIT distance="100" swimtime="00:02:39.03" />
                    <SPLIT distance="150" swimtime="00:03:58.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" status="DNS" swimtime="00:00:00.00" resultid="43535" heatid="45097" lane="2" entrytime="00:01:20.16" entrycourse="LCM" />
                <RESULT eventid="2637" points="120" swimtime="00:02:25.78" resultid="43536" heatid="44951" lane="5" entrytime="00:02:26.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" status="DNS" swimtime="00:00:00.00" resultid="43537" heatid="45117" lane="4" entrytime="00:02:51.07" entrycourse="LCM" />
                <RESULT eventid="2430" status="DNS" swimtime="00:00:00.00" resultid="43538" heatid="45066" lane="7" entrytime="00:01:03.94" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Teresa Sofia" lastname="Bento" birthdate="1974-04-13" gender="F" nation="POR" license="208407" swrid="5326683" athleteid="43209">
              <RESULTS>
                <RESULT eventid="1060" points="138" swimtime="00:18:41.86" resultid="43210" heatid="45074" lane="4" entrytime="00:18:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:02.11" />
                    <SPLIT distance="200" swimtime="00:04:17.77" />
                    <SPLIT distance="300" swimtime="00:06:39.11" />
                    <SPLIT distance="400" swimtime="00:09:08.93" />
                    <SPLIT distance="500" swimtime="00:11:38.41" />
                    <SPLIT distance="600" swimtime="00:14:03.69" />
                    <SPLIT distance="700" swimtime="00:16:31.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2173" points="198" swimtime="00:04:52.88" resultid="43211" heatid="45087" lane="8" entrytime="00:04:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.40" />
                    <SPLIT distance="100" swimtime="00:02:17.07" />
                    <SPLIT distance="150" swimtime="00:03:36.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Sofia" lastname="Silva" birthdate="1978-06-21" gender="F" nation="POR" license="206942" swrid="5277942" athleteid="43524">
              <RESULTS>
                <RESULT eventid="1060" points="506" swimtime="00:12:17.53" resultid="43525" heatid="45078" lane="1" entrytime="00:12:13.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.47" />
                    <SPLIT distance="200" swimtime="00:02:59.51" />
                    <SPLIT distance="300" swimtime="00:04:32.90" />
                    <SPLIT distance="400" swimtime="00:06:06.14" />
                    <SPLIT distance="500" swimtime="00:07:38.96" />
                    <SPLIT distance="600" swimtime="00:09:12.06" />
                    <SPLIT distance="700" swimtime="00:10:45.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2173" status="DNS" swimtime="00:00:00.00" resultid="43526" heatid="45089" lane="6" entrytime="00:03:19.69" entrycourse="LCM" />
                <RESULT eventid="2278" points="493" swimtime="00:02:46.55" resultid="43527" heatid="44904" lane="2" entrytime="00:03:02.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:20.40" />
                    <SPLIT distance="150" swimtime="00:02:03.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" status="DNS" swimtime="00:00:00.00" resultid="43528" heatid="44974" lane="8" entrytime="00:03:02.90" entrycourse="LCM" />
                <RESULT eventid="2460" status="DNS" swimtime="00:00:00.00" resultid="43529" heatid="45122" lane="4" entrytime="00:01:34.51" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antero Silva" lastname="Sousa" birthdate="1943-10-16" gender="M" nation="POR" license="205243" swrid="5231633" athleteid="43539">
              <RESULTS>
                <RESULT eventid="2622" points="323" reactiontime="+135" swimtime="00:04:57.26" resultid="43540" heatid="44873" lane="1" entrytime="00:04:54.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.61" />
                    <SPLIT distance="100" swimtime="00:02:23.40" />
                    <SPLIT distance="150" swimtime="00:03:41.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="351" reactiontime="+111" swimtime="00:00:56.09" resultid="43541" heatid="44939" lane="6" entrytime="00:00:55.95" entrycourse="LCM" />
                <RESULT eventid="2445" points="300" reactiontime="+127" swimtime="00:02:14.24" resultid="43542" heatid="44991" lane="1" entrytime="00:02:15.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="204" reactiontime="+106" swimtime="00:01:03.22" resultid="43543" heatid="45014" lane="5" entrytime="00:01:02.77" entrycourse="LCM" />
                <RESULT eventid="2652" points="150" reactiontime="+123" swimtime="00:00:58.68" resultid="43544" heatid="45033" lane="2" entrytime="00:00:56.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Americo Pedro" lastname="Goncalves" birthdate="1971-05-19" gender="M" nation="POR" license="121758" swrid="4703094" athleteid="43313">
              <RESULTS>
                <RESULT eventid="2537" points="700" reactiontime="+71" swimtime="00:01:14.16" resultid="43314" heatid="44888" lane="2" entrytime="00:01:14.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="724" reactiontime="+82" swimtime="00:00:30.77" resultid="43315" heatid="44899" lane="8" entrytime="00:00:30.98" entrycourse="LCM" />
                <RESULT eventid="2507" points="673" reactiontime="+90" swimtime="00:02:25.18" resultid="43316" heatid="45096" lane="8" entrytime="00:02:16.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                    <SPLIT distance="100" swimtime="00:01:11.57" />
                    <SPLIT distance="150" swimtime="00:01:49.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexia Alves" lastname="Fernandes" birthdate="1996-10-31" gender="F" nation="POR" license="201754" athleteid="43293">
              <RESULTS>
                <RESULT eventid="1060" points="366" swimtime="00:12:52.28" resultid="43294" heatid="45077" lane="2" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.77" />
                    <SPLIT distance="200" swimtime="00:03:03.82" />
                    <SPLIT distance="300" swimtime="00:04:41.20" />
                    <SPLIT distance="400" swimtime="00:06:20.18" />
                    <SPLIT distance="500" swimtime="00:07:59.14" />
                    <SPLIT distance="600" swimtime="00:09:37.68" />
                    <SPLIT distance="700" swimtime="00:11:16.36" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="708 - Não efectuou o ciclo completo de braçada seguida de pernada - SW 7.2" eventid="2173" status="DSQ" swimtime="00:03:43.33" resultid="43295" heatid="45088" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.01" />
                    <SPLIT distance="100" swimtime="00:01:46.76" />
                    <SPLIT distance="150" swimtime="00:02:44.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2203" points="261" reactiontime="+85" swimtime="00:01:44.04" resultid="43296" heatid="44881" lane="2" entrytime="00:01:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2338" points="255" reactiontime="+92" swimtime="00:00:43.83" resultid="43297" heatid="44889" lane="4" entrytime="00:00:55.00" />
                <RESULT eventid="2400" points="294" reactiontime="+94" swimtime="00:07:30.95" resultid="43298" heatid="45064" lane="7" entrytime="00:07:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.11" />
                    <SPLIT distance="100" swimtime="00:01:47.30" />
                    <SPLIT distance="150" swimtime="00:02:51.52" />
                    <SPLIT distance="200" swimtime="00:03:52.01" />
                    <SPLIT distance="250" swimtime="00:04:51.96" />
                    <SPLIT distance="300" swimtime="00:05:52.80" />
                    <SPLIT distance="350" swimtime="00:06:44.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jorge Manuel" lastname="Monteiro" birthdate="1967-11-28" gender="M" nation="POR" license="202134" swrid="5197050" athleteid="43384">
              <RESULTS>
                <RESULT eventid="2323" points="702" reactiontime="+78" swimtime="00:01:11.63" resultid="43385" heatid="44928" lane="4" entrytime="00:01:09.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="785" reactiontime="+77" swimtime="00:01:01.63" resultid="43386" heatid="45115" lane="1" entrytime="00:01:00.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="702" reactiontime="+93" swimtime="00:00:33.48" resultid="43387" heatid="45020" lane="5" entrytime="00:00:33.89" entrycourse="LCM" />
                <RESULT eventid="2652" points="749" reactiontime="+76" swimtime="00:00:27.65" resultid="43388" heatid="45047" lane="2" entrytime="00:00:26.88" entrycourse="LCM" />
                <RESULT eventid="2682" points="859" reactiontime="+74" swimtime="00:00:29.07" resultid="43389" heatid="44900" lane="2" entrytime="00:00:29.33" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Fonseca" lastname="Oliveira" birthdate="1974-06-13" gender="M" nation="POR" license="207947" swrid="5304477" athleteid="43416">
              <RESULTS>
                <RESULT eventid="1058" points="308" swimtime="00:13:04.36" resultid="43417" heatid="45082" lane="5" entrytime="00:13:12.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.61" />
                    <SPLIT distance="200" swimtime="00:03:07.12" />
                    <SPLIT distance="300" swimtime="00:04:43.57" />
                    <SPLIT distance="400" swimtime="00:06:22.81" />
                    <SPLIT distance="500" swimtime="00:08:04.46" />
                    <SPLIT distance="600" swimtime="00:09:44.64" />
                    <SPLIT distance="700" swimtime="00:11:27.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2537" points="206" reactiontime="+71" swimtime="00:01:44.71" resultid="43418" heatid="44886" lane="1" entrytime="00:01:37.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="227" reactiontime="+88" swimtime="00:03:42.40" resultid="43419" heatid="44918" lane="2" entrytime="00:03:46.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.90" />
                    <SPLIT distance="100" swimtime="00:01:52.27" />
                    <SPLIT distance="150" swimtime="00:02:47.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="349" reactiontime="+88" swimtime="00:01:19.26" resultid="43420" heatid="45108" lane="8" entrytime="00:01:20.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" points="207" reactiontime="+111" swimtime="00:03:55.21" resultid="43421" heatid="45029" lane="8" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.78" />
                    <SPLIT distance="100" swimtime="00:01:56.34" />
                    <SPLIT distance="150" swimtime="00:02:58.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filipa Margarida" lastname="Ferreira" birthdate="1969-03-21" gender="F" nation="POR" license="127852" swrid="4905769" athleteid="43299">
              <RESULTS>
                <RESULT eventid="2338" points="533" reactiontime="+104" swimtime="00:00:37.28" resultid="43300" heatid="44892" lane="8" entrytime="00:00:35.78" entrycourse="LCM" />
                <RESULT eventid="2607" points="554" reactiontime="+108" swimtime="00:00:44.69" resultid="43301" heatid="45101" lane="8" entrytime="00:00:48.13" entrycourse="LCM" />
                <RESULT eventid="2637" points="596" reactiontime="+106" swimtime="00:01:15.18" resultid="43302" heatid="44956" lane="1" entrytime="00:01:16.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="571" reactiontime="+70" swimtime="00:00:41.41" resultid="43303" heatid="45026" lane="6" entrytime="00:00:41.09" entrycourse="LCM" />
                <RESULT eventid="2430" points="629" reactiontime="+98" swimtime="00:00:33.15" resultid="43304" heatid="45072" lane="8" entrytime="00:00:32.05" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Giraldo" lastname="Wernicke" birthdate="1960-12-01" gender="F" nation="POR" license="210543" swrid="5367930" athleteid="43568">
              <RESULTS>
                <RESULT eventid="1060" status="DNS" swimtime="00:00:00.00" resultid="43569" heatid="45075" lane="4" entrytime="00:15:53.96" entrycourse="LCM" />
                <RESULT eventid="2203" status="DNS" swimtime="00:00:00.00" resultid="43570" heatid="44880" lane="2" entrytime="00:02:13.28" entrycourse="LCM" />
                <RESULT eventid="2278" status="DNS" swimtime="00:00:00.00" resultid="43571" heatid="44902" lane="3" entrytime="00:03:40.17" entrycourse="LCM" />
                <RESULT eventid="2492" status="DNS" swimtime="00:00:00.00" resultid="43572" heatid="45009" lane="5" entrytime="00:07:45.80" entrycourse="LCM" />
                <RESULT eventid="2430" status="DNS" swimtime="00:00:00.00" resultid="43573" heatid="45067" lane="4" entrytime="00:00:42.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Miguel" lastname="Loureiro" birthdate="1968-11-03" gender="M" nation="POR" license="205536" swrid="5277941" athleteid="43349">
              <RESULTS>
                <RESULT eventid="1058" points="190" swimtime="00:15:58.27" resultid="43350" heatid="45080" lane="2" entrytime="00:16:55.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.30" />
                    <SPLIT distance="200" swimtime="00:03:48.00" />
                    <SPLIT distance="300" swimtime="00:05:47.80" />
                    <SPLIT distance="400" swimtime="00:07:48.43" />
                    <SPLIT distance="500" swimtime="00:09:50.53" />
                    <SPLIT distance="600" swimtime="00:11:52.76" />
                    <SPLIT distance="700" swimtime="00:13:56.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="230" reactiontime="+111" swimtime="00:01:32.75" resultid="43351" heatid="45104" lane="5" entrytime="00:01:41.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="193" reactiontime="+117" swimtime="00:07:42.32" resultid="43352" heatid="45125" lane="8" entrytime="00:08:15.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.84" />
                    <SPLIT distance="100" swimtime="00:01:41.55" />
                    <SPLIT distance="150" swimtime="00:02:39.83" />
                    <SPLIT distance="200" swimtime="00:03:39.37" />
                    <SPLIT distance="250" swimtime="00:04:40.44" />
                    <SPLIT distance="300" swimtime="00:05:41.28" />
                    <SPLIT distance="350" swimtime="00:06:42.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Rosa" lastname="Palhares" birthdate="1965-06-22" gender="F" nation="POR" license="201379" swrid="5171502" athleteid="43422">
              <RESULTS>
                <RESULT eventid="2607" status="DNS" swimtime="00:00:00.00" resultid="43423" heatid="45100" lane="3" entrytime="00:00:49.02" entrycourse="LCM" />
                <RESULT eventid="2637" status="DNS" swimtime="00:00:00.00" resultid="43424" heatid="44953" lane="5" entrytime="00:01:37.00" entrycourse="LCM" />
                <RESULT eventid="2460" status="DNS" swimtime="00:00:00.00" resultid="43425" heatid="45120" lane="8" entrytime="00:01:56.75" entrycourse="LCM" />
                <RESULT eventid="2492" status="DNS" swimtime="00:00:00.00" resultid="43426" heatid="45009" lane="1" entrytime="00:08:07.45" entrycourse="LCM" />
                <RESULT eventid="2522" status="DNS" swimtime="00:00:00.00" resultid="43427" heatid="45024" lane="1" entrytime="00:00:54.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Castro" lastname="Rocha" birthdate="1995-06-07" gender="M" nation="POR" license="212348" swrid="5424187" athleteid="43482">
              <RESULTS>
                <RESULT eventid="1058" points="117" swimtime="00:17:43.52" resultid="43483" heatid="45080" lane="7" entrytime="00:17:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.14" />
                    <SPLIT distance="200" swimtime="00:04:00.14" />
                    <SPLIT distance="300" swimtime="00:06:15.55" />
                    <SPLIT distance="400" swimtime="00:08:33.00" />
                    <SPLIT distance="500" swimtime="00:10:49.88" />
                    <SPLIT distance="600" swimtime="00:13:08.08" />
                    <SPLIT distance="700" swimtime="00:15:26.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2622" points="194" reactiontime="+149" swimtime="00:04:09.77" resultid="43484" heatid="44874" lane="1" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.07" />
                    <SPLIT distance="100" swimtime="00:02:00.34" />
                    <SPLIT distance="150" swimtime="00:03:05.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="118" reactiontime="+130" swimtime="00:03:54.33" resultid="43485" heatid="45090" lane="6" entrytime="00:04:11.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.02" />
                    <SPLIT distance="100" swimtime="00:01:49.34" />
                    <SPLIT distance="150" swimtime="00:02:50.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="120" reactiontime="+130" swimtime="00:08:27.45" resultid="43486" heatid="45124" lane="3" entrytime="00:08:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.58" />
                    <SPLIT distance="100" swimtime="00:01:51.80" />
                    <SPLIT distance="150" swimtime="00:02:55.26" />
                    <SPLIT distance="200" swimtime="00:04:02.86" />
                    <SPLIT distance="250" swimtime="00:05:08.36" />
                    <SPLIT distance="300" swimtime="00:06:16.94" />
                    <SPLIT distance="350" swimtime="00:07:24.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sergio Manuel" lastname="Neves" birthdate="1982-10-02" gender="M" nation="POR" license="204875" swrid="5215134" athleteid="43405">
              <RESULTS>
                <RESULT eventid="2622" points="205" reactiontime="+101" swimtime="00:04:16.53" resultid="43406" heatid="44873" lane="4" entrytime="00:04:19.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.56" />
                    <SPLIT distance="100" swimtime="00:02:09.84" />
                    <SPLIT distance="150" swimtime="00:03:16.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="146" reactiontime="+96" swimtime="00:03:39.67" resultid="43407" heatid="45090" lane="5" entrytime="00:03:49.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.47" />
                    <SPLIT distance="100" swimtime="00:01:47.78" />
                    <SPLIT distance="150" swimtime="00:02:46.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="148" reactiontime="+89" swimtime="00:04:11.68" resultid="43408" heatid="44917" lane="3" entrytime="00:04:07.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.54" />
                    <SPLIT distance="100" swimtime="00:02:08.66" />
                    <SPLIT distance="150" swimtime="00:03:13.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="169" reactiontime="+102" swimtime="00:03:58.55" resultid="43409" heatid="44976" lane="1" entrytime="00:04:02.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.79" />
                    <SPLIT distance="100" swimtime="00:02:02.93" />
                    <SPLIT distance="150" swimtime="00:03:07.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="124" reactiontime="+104" swimtime="00:08:34.10" resultid="43410" heatid="45125" lane="7" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.32" />
                    <SPLIT distance="100" swimtime="00:01:57.47" />
                    <SPLIT distance="150" swimtime="00:03:07.41" />
                    <SPLIT distance="200" swimtime="00:04:18.75" />
                    <SPLIT distance="250" swimtime="00:05:28.45" />
                    <SPLIT distance="300" swimtime="00:06:35.87" />
                    <SPLIT distance="350" swimtime="00:07:40.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Luis" lastname="Roseira" birthdate="1955-02-27" gender="M" nation="POR" license="142204" swrid="5119322" athleteid="43492">
              <RESULTS>
                <RESULT eventid="2622" points="164" reactiontime="+116" swimtime="00:05:42.21" resultid="43493" heatid="44873" lane="8" entrytime="00:05:03.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.17" />
                    <SPLIT distance="100" swimtime="00:02:48.03" />
                    <SPLIT distance="150" swimtime="00:04:17.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="65" reactiontime="+130" swimtime="00:01:15.72" resultid="43494" heatid="44893" lane="1" entrytime="00:01:09.52" entrycourse="LCM" />
                <RESULT eventid="2188" points="181" reactiontime="+129" swimtime="00:01:00.92" resultid="43495" heatid="44939" lane="7" entrytime="00:00:59.73" entrycourse="LCM" />
                <RESULT eventid="2445" points="169" reactiontime="+122" swimtime="00:02:28.74" resultid="43496" heatid="44991" lane="6" entrytime="00:02:14.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="185" reactiontime="+116" swimtime="00:00:49.73" resultid="43497" heatid="45034" lane="8" entrytime="00:00:46.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Luis" lastname="Morgado" birthdate="1954-03-14" gender="M" nation="POR" license="124934" swrid="4005115" athleteid="43390">
              <RESULTS>
                <RESULT eventid="2188" points="239" reactiontime="+109" swimtime="00:00:55.56" resultid="43391" heatid="44941" lane="6" entrytime="00:00:48.65" entrycourse="LCM" />
                <RESULT eventid="2415" points="299" reactiontime="+108" swimtime="00:01:33.81" resultid="43392" heatid="45106" lane="5" entrytime="00:01:26.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="288" reactiontime="+114" swimtime="00:02:04.70" resultid="43393" heatid="44992" lane="7" entrytime="00:01:58.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="227" reactiontime="+85" swimtime="00:00:54.89" resultid="43394" heatid="45015" lane="2" entrytime="00:00:56.44" entrycourse="LCM" />
                <RESULT eventid="2652" points="367" reactiontime="+100" swimtime="00:00:39.62" resultid="43395" heatid="45036" lane="6" entrytime="00:00:37.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui David" lastname="Castro" birthdate="1970-01-01" gender="M" nation="POR" license="214263" athleteid="43256">
              <RESULTS>
                <RESULT eventid="2323" points="574" reactiontime="+96" swimtime="00:01:16.60" resultid="43257" heatid="44928" lane="7" entrytime="00:01:13.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="619" reactiontime="+89" swimtime="00:01:06.70" resultid="43258" heatid="45113" lane="2" entrytime="00:01:04.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="673" reactiontime="+95" swimtime="00:00:31.53" resultid="43259" heatid="44898" lane="4" entrytime="00:00:31.00" />
                <RESULT eventid="2652" points="639" reactiontime="+95" swimtime="00:00:29.15" resultid="43260" heatid="45046" lane="6" entrytime="00:00:27.50" />
                <RESULT eventid="2248" points="478" reactiontime="+100" swimtime="00:06:45.71" resultid="43261" heatid="45061" lane="1" entrytime="00:06:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                    <SPLIT distance="100" swimtime="00:01:25.19" />
                    <SPLIT distance="150" swimtime="00:02:26.12" />
                    <SPLIT distance="200" swimtime="00:03:24.32" />
                    <SPLIT distance="250" swimtime="00:04:24.68" />
                    <SPLIT distance="300" swimtime="00:05:22.71" />
                    <SPLIT distance="350" swimtime="00:06:06.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paula Alexandra" lastname="Palhares" birthdate="1966-09-27" gender="F" nation="POR" license="212331" swrid="5424178" athleteid="43434">
              <RESULTS>
                <RESULT eventid="2203" points="556" reactiontime="+80" swimtime="00:01:34.98" resultid="43435" heatid="44883" lane="1" entrytime="00:01:29.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2278" points="376" reactiontime="+109" swimtime="00:03:13.56" resultid="43436" heatid="44904" lane="4" entrytime="00:02:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                    <SPLIT distance="100" swimtime="00:01:28.71" />
                    <SPLIT distance="150" swimtime="00:02:20.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2308" points="487" reactiontime="+89" swimtime="00:03:32.16" resultid="43437" heatid="44915" lane="8" entrytime="00:03:15.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.28" />
                    <SPLIT distance="100" swimtime="00:01:43.78" />
                    <SPLIT distance="150" swimtime="00:02:38.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="578" reactiontime="+80" swimtime="00:00:42.90" resultid="43438" heatid="45026" lane="3" entrytime="00:00:40.96" entrycourse="SCM" />
                <RESULT eventid="2430" points="526" reactiontime="+100" swimtime="00:00:36.67" resultid="43439" heatid="45070" lane="2" entrytime="00:00:35.57" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Lopes" lastname="Santos" birthdate="1959-03-21" gender="M" nation="POR" license="124875" swrid="4005259" athleteid="43512">
              <RESULTS>
                <RESULT eventid="2682" points="602" reactiontime="+86" swimtime="00:00:34.47" resultid="43513" heatid="44896" lane="5" entrytime="00:00:35.70" entrycourse="SCM" />
                <RESULT eventid="2188" status="DNS" swimtime="00:00:00.00" resultid="43514" heatid="44946" lane="2" entrytime="00:00:41.01" entrycourse="LCM" />
                <RESULT eventid="2415" points="608" reactiontime="+91" swimtime="00:01:12.03" resultid="43515" heatid="45110" lane="6" entrytime="00:01:11.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="541" reactiontime="+63" swimtime="00:00:40.38" resultid="43516" heatid="45019" lane="8" entrytime="00:00:40.42" entrycourse="LCM" />
                <RESULT eventid="2652" points="694" reactiontime="+93" swimtime="00:00:30.86" resultid="43517" heatid="45042" lane="8" entrytime="00:00:30.41" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ines Maria" lastname="Rothes" birthdate="1973-12-16" gender="F" nation="POR" license="124731" swrid="4564410" athleteid="43498">
              <RESULTS>
                <RESULT eventid="1060" points="432" swimtime="00:12:47.80" resultid="43499" heatid="45078" lane="3" entrytime="00:11:20.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.84" />
                    <SPLIT distance="200" swimtime="00:03:00.87" />
                    <SPLIT distance="300" swimtime="00:04:37.76" />
                    <SPLIT distance="400" swimtime="00:06:06.36" />
                    <SPLIT distance="500" swimtime="00:07:54.61" />
                    <SPLIT distance="600" swimtime="00:09:33.02" />
                    <SPLIT distance="700" swimtime="00:11:11.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="450" swimtime="00:06:10.99" resultid="43500" heatid="45013" lane="3" entrytime="00:05:25.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.30" />
                    <SPLIT distance="100" swimtime="00:01:24.53" />
                    <SPLIT distance="150" swimtime="00:02:10.66" />
                    <SPLIT distance="200" swimtime="00:02:58.60" />
                    <SPLIT distance="250" swimtime="00:03:47.40" />
                    <SPLIT distance="300" swimtime="00:04:35.51" />
                    <SPLIT distance="350" swimtime="00:05:23.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Nuno" lastname="Goncalves" birthdate="1972-05-25" gender="M" nation="POR" license="205032" swrid="5227009" athleteid="43323">
              <RESULTS>
                <RESULT eventid="1058" points="187" swimtime="00:15:25.65" resultid="43324" heatid="45081" lane="8" entrytime="00:15:33.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.03" />
                    <SPLIT distance="200" swimtime="00:03:46.02" />
                    <SPLIT distance="300" swimtime="00:05:45.01" />
                    <SPLIT distance="400" swimtime="00:07:43.36" />
                    <SPLIT distance="500" swimtime="00:09:42.99" />
                    <SPLIT distance="600" swimtime="00:11:41.68" />
                    <SPLIT distance="700" swimtime="00:13:37.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2537" points="82" reactiontime="+94" swimtime="00:02:21.98" resultid="43325" heatid="44884" lane="3" entrytime="00:02:16.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Margarida Maria" lastname="Ribeiro" birthdate="1964-06-04" gender="F" nation="POR" license="131782" swrid="5036828" athleteid="43476">
              <RESULTS>
                <RESULT eventid="2308" points="119" reactiontime="+118" swimtime="00:05:39.35" resultid="43477" heatid="44913" lane="1" entrytime="00:05:14.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:24.57" />
                    <SPLIT distance="100" swimtime="00:02:50.90" />
                    <SPLIT distance="150" swimtime="00:04:16.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="147" reactiontime="+121" swimtime="00:02:00.64" resultid="43478" heatid="44952" lane="7" entrytime="00:02:07.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="96" reactiontime="+132" swimtime="00:05:46.47" resultid="43479" heatid="44971" lane="7" entrytime="00:05:08.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:23.04" />
                    <SPLIT distance="100" swimtime="00:03:01.22" />
                    <SPLIT distance="150" swimtime="00:04:31.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="111" reactiontime="+136" swimtime="00:01:14.30" resultid="43480" heatid="45023" lane="2" entrytime="00:01:06.83" entrycourse="LCM" />
                <RESULT eventid="2430" points="185" reactiontime="+126" swimtime="00:00:51.88" resultid="43481" heatid="45067" lane="8" entrytime="00:00:49.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leandro Filipe" lastname="Sousa" birthdate="1972-01-13" gender="M" nation="POR" license="204933" swrid="5220452" athleteid="43545">
              <RESULTS>
                <RESULT eventid="2682" points="464" reactiontime="+90" swimtime="00:00:34.30" resultid="43546" heatid="44897" lane="5" entrytime="00:00:33.22" entrycourse="LCM" />
                <RESULT eventid="2507" points="430" reactiontime="+92" swimtime="00:02:38.08" resultid="43547" heatid="45094" lane="4" entrytime="00:02:28.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="100" swimtime="00:01:15.37" />
                    <SPLIT distance="150" swimtime="00:01:57.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2323" points="365" reactiontime="+99" swimtime="00:01:24.51" resultid="43548" heatid="44927" lane="2" entrytime="00:01:21.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="620" reactiontime="+84" swimtime="00:01:05.47" resultid="43549" heatid="45112" lane="6" entrytime="00:01:05.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carla Susana" lastname="Avelans" birthdate="1975-05-10" gender="F" nation="POR" license="130741" swrid="5003421" athleteid="43194">
              <RESULTS>
                <RESULT eventid="2173" points="421" swimtime="00:03:48.06" resultid="43195" heatid="45088" lane="4" entrytime="00:03:42.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.88" />
                    <SPLIT distance="100" swimtime="00:01:49.98" />
                    <SPLIT distance="150" swimtime="00:02:49.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2203" points="241" reactiontime="+112" swimtime="00:01:53.00" resultid="43196" heatid="44881" lane="3" entrytime="00:01:49.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2308" points="299" reactiontime="+104" swimtime="00:03:57.93" resultid="43197" heatid="44914" lane="2" entrytime="00:03:50.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.49" />
                    <SPLIT distance="100" swimtime="00:01:56.65" />
                    <SPLIT distance="150" swimtime="00:02:56.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="437" reactiontime="+105" swimtime="00:01:45.52" resultid="43198" heatid="45121" lane="5" entrytime="00:01:41.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" status="DNS" swimtime="00:00:00.00" resultid="43199" heatid="45009" lane="7" entrytime="00:07:54.57" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Pedro" lastname="Santana" birthdate="1966-09-05" gender="M" nation="POR" license="124877" swrid="4005248" athleteid="43507">
              <RESULTS>
                <RESULT eventid="2682" status="DNS" swimtime="00:00:00.00" resultid="43508" heatid="44898" lane="5" entrytime="00:00:31.05" entrycourse="LCM" />
                <RESULT eventid="2188" status="DNS" swimtime="00:00:00.00" resultid="43509" heatid="44949" lane="3" entrytime="00:00:35.27" entrycourse="LCM" />
                <RESULT eventid="2293" status="DNS" swimtime="00:00:00.00" resultid="43510" heatid="45020" lane="3" entrytime="00:00:34.25" entrycourse="LCM" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="43511" heatid="45045" lane="2" entrytime="00:00:28.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lilia Dulce" lastname="Costa" birthdate="1981-12-08" gender="F" nation="POR" license="132418" swrid="5068111" athleteid="43271">
              <RESULTS>
                <RESULT eventid="2492" points="358" reactiontime="+90" swimtime="00:06:38.06" resultid="43272" heatid="45012" lane="3" entrytime="00:06:16.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.85" />
                    <SPLIT distance="100" swimtime="00:01:25.49" />
                    <SPLIT distance="150" swimtime="00:02:16.18" />
                    <SPLIT distance="200" swimtime="00:03:08.59" />
                    <SPLIT distance="250" swimtime="00:04:01.26" />
                    <SPLIT distance="300" swimtime="00:04:55.40" />
                    <SPLIT distance="350" swimtime="00:05:46.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="368" reactiontime="+72" swimtime="00:00:44.19" resultid="43273" heatid="45026" lane="7" entrytime="00:00:41.32" entrycourse="SCM" />
                <RESULT eventid="2430" points="438" reactiontime="+84" swimtime="00:00:36.12" resultid="43274" heatid="45069" lane="3" entrytime="00:00:37.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Sofia" lastname="Uhlfelder" birthdate="1983-10-05" gender="F" nation="POR" license="200872" swrid="5159395" athleteid="43556">
              <RESULTS>
                <RESULT eventid="2552" points="171" reactiontime="+125" swimtime="00:01:59.87" resultid="43557" heatid="44923" lane="1" entrytime="00:02:01.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="165" reactiontime="+119" swimtime="00:00:59.45" resultid="43558" heatid="45098" lane="7" entrytime="00:00:59.63" entrycourse="SCM" />
                <RESULT eventid="2637" points="241" reactiontime="+113" swimtime="00:01:35.52" resultid="43559" heatid="44953" lane="2" entrytime="00:01:45.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="236" reactiontime="+110" swimtime="00:04:01.07" resultid="43560" heatid="44972" lane="8" entrytime="00:04:05.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.00" />
                    <SPLIT distance="100" swimtime="00:01:54.10" />
                    <SPLIT distance="150" swimtime="00:03:05.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="192" reactiontime="+124" swimtime="00:02:05.67" resultid="43561" heatid="45119" lane="1" entrytime="00:02:05.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos Guimaraes" lastname="Goncalves" birthdate="1970-11-22" gender="M" nation="POR" license="123664" swrid="4763854" athleteid="43317">
              <RESULTS>
                <RESULT eventid="2248" points="615" reactiontime="+92" swimtime="00:06:13.16" resultid="43318" heatid="45061" lane="5" entrytime="00:06:02.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                    <SPLIT distance="100" swimtime="00:01:15.61" />
                    <SPLIT distance="150" swimtime="00:02:04.53" />
                    <SPLIT distance="200" swimtime="00:02:53.74" />
                    <SPLIT distance="250" swimtime="00:03:50.57" />
                    <SPLIT distance="300" swimtime="00:04:47.63" />
                    <SPLIT distance="350" swimtime="00:05:30.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1058" points="501" swimtime="00:11:33.71" resultid="43319" heatid="45085" lane="3" entrytime="00:10:27.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.11" />
                    <SPLIT distance="200" swimtime="00:02:43.22" />
                    <SPLIT distance="300" swimtime="00:04:08.44" />
                    <SPLIT distance="400" swimtime="00:05:36.27" />
                    <SPLIT distance="500" swimtime="00:07:05.14" />
                    <SPLIT distance="600" swimtime="00:08:35.12" />
                    <SPLIT distance="700" swimtime="00:10:05.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2622" points="517" reactiontime="+101" swimtime="00:03:19.40" resultid="43320" heatid="44877" lane="5" entrytime="00:03:18.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.96" />
                    <SPLIT distance="100" swimtime="00:01:38.03" />
                    <SPLIT distance="150" swimtime="00:02:28.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2537" points="551" reactiontime="+88" swimtime="00:01:20.32" resultid="43321" heatid="44888" lane="7" entrytime="00:01:14.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="633" reactiontime="+87" swimtime="00:02:28.16" resultid="43322" heatid="45095" lane="5" entrytime="00:02:19.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                    <SPLIT distance="100" swimtime="00:01:11.37" />
                    <SPLIT distance="150" swimtime="00:01:50.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Alberto" lastname="Mendes" birthdate="1975-10-11" gender="M" nation="POR" license="202097" swrid="5197049" athleteid="43375">
              <RESULTS>
                <RESULT eventid="1058" points="351" swimtime="00:12:31.11" resultid="43376" heatid="45083" lane="8" entrytime="00:13:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.08" />
                    <SPLIT distance="200" swimtime="00:02:55.15" />
                    <SPLIT distance="300" swimtime="00:04:30.02" />
                    <SPLIT distance="400" swimtime="00:06:05.88" />
                    <SPLIT distance="500" swimtime="00:07:42.55" />
                    <SPLIT distance="600" swimtime="00:09:19.64" />
                    <SPLIT distance="700" swimtime="00:10:56.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2537" points="302" reactiontime="+78" swimtime="00:01:32.13" resultid="43377" heatid="44887" lane="1" entrytime="00:01:29.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="467" reactiontime="+98" swimtime="00:01:11.98" resultid="43378" heatid="45109" lane="4" entrytime="00:01:13.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="394" swimtime="00:00:39.24" resultid="43379" heatid="45018" lane="6" entrytime="00:00:42.93" entrycourse="LCM" />
                <RESULT eventid="2652" points="451" reactiontime="+95" swimtime="00:00:32.43" resultid="43380" heatid="45040" lane="1" entrytime="00:00:32.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Miguel" lastname="Barroso" birthdate="1962-05-19" gender="M" nation="POR" license="208445" swrid="5326682" athleteid="43203">
              <RESULTS>
                <RESULT eventid="2622" points="644" reactiontime="+88" swimtime="00:03:09.27" resultid="43204" heatid="44878" lane="1" entrytime="00:03:15.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.79" />
                    <SPLIT distance="100" swimtime="00:01:31.88" />
                    <SPLIT distance="150" swimtime="00:02:20.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="557" reactiontime="+85" swimtime="00:02:37.44" resultid="43205" heatid="45093" lane="5" entrytime="00:02:42.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                    <SPLIT distance="100" swimtime="00:01:13.07" />
                    <SPLIT distance="150" swimtime="00:01:54.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="591" reactiontime="+75" swimtime="00:00:36.99" resultid="43206" heatid="44948" lane="2" entrytime="00:00:37.98" entrycourse="LCM" />
                <RESULT eventid="2445" points="674" reactiontime="+86" swimtime="00:01:22.82" resultid="43207" heatid="44998" lane="7" entrytime="00:01:24.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" status="DNS" swimtime="00:00:00.00" resultid="43208" heatid="45127" lane="7" entrytime="00:06:43.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Gunther" lastname="Amaral" birthdate="1969-07-19" gender="M" nation="POR" license="209669" swrid="5344157" athleteid="43183">
              <RESULTS>
                <RESULT eventid="2622" points="363" reactiontime="+92" swimtime="00:03:44.25" resultid="43184" heatid="44877" lane="8" entrytime="00:03:24.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.07" />
                    <SPLIT distance="100" swimtime="00:01:43.40" />
                    <SPLIT distance="150" swimtime="00:02:42.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="333" reactiontime="+89" swimtime="00:00:44.90" resultid="43185" heatid="44943" lane="5" entrytime="00:00:44.50" entrycourse="LCM" />
                <RESULT eventid="2415" points="275" reactiontime="+87" swimtime="00:01:27.43" resultid="43186" heatid="45105" lane="3" entrytime="00:01:31.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="364" reactiontime="+96" swimtime="00:01:41.51" resultid="43187" heatid="44993" lane="4" entrytime="00:01:44.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta Sofia" lastname="Oliveira" birthdate="1983-12-13" gender="F" nation="POR" license="128880" swrid="4938968" athleteid="43411">
              <RESULTS>
                <RESULT eventid="2637" points="623" reactiontime="+88" swimtime="00:01:09.61" resultid="43412" heatid="44957" lane="1" entrytime="00:01:10.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="507" reactiontime="+74" swimtime="00:03:07.02" resultid="43413" heatid="44973" lane="4" entrytime="00:03:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                    <SPLIT distance="100" swimtime="00:01:25.21" />
                    <SPLIT distance="150" swimtime="00:02:23.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="541" reactiontime="+75" swimtime="00:00:39.32" resultid="43414" heatid="45027" lane="1" entrytime="00:00:38.36" entrycourse="LCM" />
                <RESULT eventid="2430" points="690" reactiontime="+79" swimtime="00:00:30.37" resultid="43415" heatid="45073" lane="6" entrytime="00:00:29.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joana Isabel" lastname="Leite" birthdate="1980-01-06" gender="F" nation="POR" license="130666" swrid="5001721" athleteid="43332">
              <RESULTS>
                <RESULT eventid="1060" points="132" swimtime="00:19:13.13" resultid="43333" heatid="45075" lane="7" entrytime="00:17:31.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:09.46" />
                    <SPLIT distance="200" swimtime="00:04:31.16" />
                    <SPLIT distance="300" swimtime="00:06:57.47" />
                    <SPLIT distance="400" swimtime="00:09:22.86" />
                    <SPLIT distance="500" swimtime="00:11:49.91" />
                    <SPLIT distance="600" swimtime="00:14:20.80" />
                    <SPLIT distance="700" swimtime="00:16:50.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2173" points="341" swimtime="00:04:03.06" resultid="43334" heatid="45088" lane="7" entrytime="00:03:57.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.11" />
                    <SPLIT distance="100" swimtime="00:01:56.71" />
                    <SPLIT distance="150" swimtime="00:03:00.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2203" points="200" reactiontime="+133" swimtime="00:01:59.73" resultid="43335" heatid="44880" lane="3" entrytime="00:02:03.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2308" points="242" reactiontime="+104" swimtime="00:04:06.83" resultid="43336" heatid="44913" lane="4" entrytime="00:04:08.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.63" />
                    <SPLIT distance="100" swimtime="00:02:01.76" />
                    <SPLIT distance="150" swimtime="00:03:04.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="148" swimtime="00:08:53.42" resultid="43337" heatid="45008" lane="4" entrytime="00:08:17.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.14" />
                    <SPLIT distance="100" swimtime="00:02:03.01" />
                    <SPLIT distance="150" swimtime="00:03:11.55" />
                    <SPLIT distance="200" swimtime="00:04:19.68" />
                    <SPLIT distance="250" swimtime="00:05:29.16" />
                    <SPLIT distance="300" swimtime="00:06:37.03" />
                    <SPLIT distance="350" swimtime="00:07:45.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filipe Miguel" lastname="Silva" birthdate="1974-09-28" gender="M" nation="POR" license="201375" swrid="5171525" athleteid="43530">
              <RESULTS>
                <RESULT eventid="2218" points="239" reactiontime="+75" swimtime="00:03:38.47" resultid="43531" heatid="44918" lane="5" entrytime="00:03:37.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.60" />
                    <SPLIT distance="100" swimtime="00:01:47.39" />
                    <SPLIT distance="150" swimtime="00:02:45.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="292" reactiontime="+85" swimtime="00:03:27.48" resultid="43532" heatid="44976" lane="4" entrytime="00:03:40.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.40" />
                    <SPLIT distance="100" swimtime="00:01:42.56" />
                    <SPLIT distance="150" swimtime="00:02:42.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Rui" lastname="Amaral" birthdate="1963-02-23" gender="M" nation="POR" license="206897" swrid="5276256" athleteid="43188">
              <RESULTS>
                <RESULT eventid="1058" points="320" swimtime="00:13:48.77" resultid="43189" heatid="45082" lane="6" entrytime="00:13:37.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:03:22.61" />
                    <SPLIT distance="300" swimtime="00:05:08.28" />
                    <SPLIT distance="400" swimtime="00:06:53.55" />
                    <SPLIT distance="500" swimtime="00:08:38.70" />
                    <SPLIT distance="600" swimtime="00:10:24.35" />
                    <SPLIT distance="700" swimtime="00:12:09.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="354" reactiontime="+123" swimtime="00:03:03.13" resultid="43190" heatid="45092" lane="7" entrytime="00:03:02.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                    <SPLIT distance="100" swimtime="00:01:28.28" />
                    <SPLIT distance="150" swimtime="00:02:17.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2323" points="158" reactiontime="+105" swimtime="00:01:59.53" resultid="43191" heatid="44926" lane="8" entrytime="00:01:55.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="384" reactiontime="+99" swimtime="00:01:22.64" resultid="43192" heatid="45107" lane="5" entrytime="00:01:21.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="338" reactiontime="+99" swimtime="00:06:36.29" resultid="43193" heatid="45127" lane="4" entrytime="00:06:29.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                    <SPLIT distance="100" swimtime="00:01:30.89" />
                    <SPLIT distance="150" swimtime="00:02:19.82" />
                    <SPLIT distance="200" swimtime="00:03:11.44" />
                    <SPLIT distance="250" swimtime="00:04:03.27" />
                    <SPLIT distance="300" swimtime="00:04:55.65" />
                    <SPLIT distance="350" swimtime="00:05:49.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Flavio Miguel" lastname="Barbara" birthdate="1995-12-11" gender="M" nation="POR" license="119741" swrid="4610210" athleteid="43200">
              <RESULTS>
                <RESULT eventid="2293" status="DNS" swimtime="00:00:00.00" resultid="43201" heatid="45021" lane="6" entrytime="00:00:33.00" />
                <RESULT eventid="2652" points="702" reactiontime="+64" swimtime="00:00:26.04" resultid="43202" heatid="45047" lane="7" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Alves" lastname="Cecilio" birthdate="1954-04-10" gender="M" nation="POR" license="100919" swrid="4403439" athleteid="43262">
              <RESULTS>
                <RESULT eventid="2622" points="516" reactiontime="+113" swimtime="00:03:53.79" resultid="43263" heatid="44875" lane="4" entrytime="00:03:38.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.46" />
                    <SPLIT distance="100" swimtime="00:01:51.65" />
                    <SPLIT distance="150" swimtime="00:02:54.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2537" points="272" reactiontime="+80" swimtime="00:01:53.80" resultid="43264" heatid="44885" lane="6" entrytime="00:01:53.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="375" reactiontime="+111" swimtime="00:00:47.84" resultid="43265" heatid="44943" lane="3" entrytime="00:00:44.71" entrycourse="LCM" />
                <RESULT eventid="2445" points="440" reactiontime="+109" swimtime="00:01:48.23" resultid="43266" heatid="44995" lane="5" entrytime="00:01:37.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="270" reactiontime="+98" swimtime="00:00:51.79" resultid="43267" heatid="45016" lane="4" entrytime="00:00:48.41" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco David" lastname="Ferreira" birthdate="1989-07-25" gender="M" nation="POR" license="121874" swrid="4574825" athleteid="43305">
              <RESULTS>
                <RESULT eventid="2415" points="498" reactiontime="+94" swimtime="00:01:04.12" resultid="43306" heatid="45111" lane="4" entrytime="00:01:06.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="473" reactiontime="+86" swimtime="00:02:48.81" resultid="43307" heatid="44981" lane="1" entrytime="00:02:45.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                    <SPLIT distance="100" swimtime="00:01:18.70" />
                    <SPLIT distance="150" swimtime="00:02:08.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1058" points="355" swimtime="00:11:29.30" resultid="43308" heatid="45084" lane="7" entrytime="00:12:00.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.51" />
                    <SPLIT distance="200" swimtime="00:02:40.94" />
                    <SPLIT distance="300" swimtime="00:04:06.96" />
                    <SPLIT distance="400" swimtime="00:05:33.44" />
                    <SPLIT distance="500" swimtime="00:07:02.00" />
                    <SPLIT distance="600" swimtime="00:08:31.51" />
                    <SPLIT distance="700" swimtime="00:10:01.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="467" reactiontime="+97" swimtime="00:05:20.15" resultid="43309" heatid="45130" lane="4" entrytime="00:05:19.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                    <SPLIT distance="100" swimtime="00:01:12.84" />
                    <SPLIT distance="150" swimtime="00:01:52.53" />
                    <SPLIT distance="200" swimtime="00:02:33.09" />
                    <SPLIT distance="250" swimtime="00:03:14.73" />
                    <SPLIT distance="300" swimtime="00:03:56.98" />
                    <SPLIT distance="350" swimtime="00:04:39.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="461" reactiontime="+98" swimtime="00:02:29.73" resultid="43310" heatid="45095" lane="7" entrytime="00:02:26.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="100" swimtime="00:01:09.54" />
                    <SPLIT distance="150" swimtime="00:01:49.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sara Cristina" lastname="Campos" birthdate="1973-06-09" gender="F" nation="POR" license="212605" swrid="5429039" athleteid="43230">
              <RESULTS>
                <RESULT eventid="2607" points="356" reactiontime="+117" swimtime="00:00:51.07" resultid="43231" heatid="45100" lane="8" entrytime="00:00:50.53" entrycourse="SCM" />
                <RESULT eventid="2460" points="373" reactiontime="+110" swimtime="00:01:51.27" resultid="43232" heatid="45119" lane="5" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Astride" lastname="Almeida" birthdate="1972-02-03" gender="F" nation="POR" license="212350" swrid="5424149" athleteid="43178">
              <RESULTS>
                <RESULT eventid="1060" points="122" swimtime="00:19:28.80" resultid="43179" heatid="45074" lane="5" entrytime="00:18:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:14.65" />
                    <SPLIT distance="200" swimtime="00:04:41.31" />
                    <SPLIT distance="300" swimtime="00:07:10.41" />
                    <SPLIT distance="400" swimtime="00:09:38.46" />
                    <SPLIT distance="500" swimtime="00:12:06.51" />
                    <SPLIT distance="600" swimtime="00:14:36.70" />
                    <SPLIT distance="700" swimtime="00:17:04.62" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="705 - Saiu na posição dorsal após a partida - SW 7.2" eventid="2173" status="DSQ" swimtime="00:04:20.75" resultid="43180" heatid="45087" lane="7" entrytime="00:04:25.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.35" />
                    <SPLIT distance="100" swimtime="00:02:12.49" />
                    <SPLIT distance="150" swimtime="00:03:18.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos Fernandes" lastname="Queiros" birthdate="1986-10-27" gender="M" nation="POR" license="118205" swrid="4123926" athleteid="43471">
              <RESULTS>
                <RESULT eventid="2507" status="DNS" swimtime="00:00:00.00" resultid="43472" heatid="45096" lane="6" entrytime="00:02:11.00" />
                <RESULT eventid="2415" points="676" reactiontime="+72" swimtime="00:00:59.20" resultid="43473" heatid="45116" lane="7" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="638" reactiontime="+74" swimtime="00:04:57.97" resultid="43474" heatid="45131" lane="6" entrytime="00:04:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.67" />
                    <SPLIT distance="100" swimtime="00:01:09.25" />
                    <SPLIT distance="150" swimtime="00:01:47.07" />
                    <SPLIT distance="200" swimtime="00:02:24.32" />
                    <SPLIT distance="250" swimtime="00:03:02.03" />
                    <SPLIT distance="300" swimtime="00:03:39.76" />
                    <SPLIT distance="350" swimtime="00:04:18.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="726" reactiontime="+68" swimtime="00:00:26.17" resultid="43475" heatid="45048" lane="7" entrytime="00:00:26.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Mota" lastname="Costa" birthdate="1971-02-21" gender="M" nation="POR" license="129079" swrid="4951635" athleteid="43281">
              <RESULTS>
                <RESULT eventid="2188" points="555" reactiontime="+86" swimtime="00:00:37.88" resultid="43282" heatid="44947" lane="8" entrytime="00:00:39.52" entrycourse="LCM" />
                <RESULT eventid="2415" points="589" reactiontime="+86" swimtime="00:01:07.83" resultid="43283" heatid="45112" lane="1" entrytime="00:01:06.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="573" reactiontime="+81" swimtime="00:01:27.24" resultid="43284" heatid="44997" lane="7" entrytime="00:01:28.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Abel" lastname="Pereira" birthdate="1973-11-12" gender="M" nation="POR" license="153155" swrid="5112981" athleteid="43444">
              <RESULTS>
                <RESULT eventid="2682" points="232" reactiontime="+118" swimtime="00:00:43.21" resultid="43445" heatid="44893" lane="4" entrytime="00:00:47.71" entrycourse="LCM" />
                <RESULT eventid="2507" points="197" reactiontime="+125" swimtime="00:03:24.95" resultid="43446" heatid="45091" lane="3" entrytime="00:03:20.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.22" />
                    <SPLIT distance="100" swimtime="00:01:39.12" />
                    <SPLIT distance="150" swimtime="00:02:34.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="137" reactiontime="+132" swimtime="00:04:22.61" resultid="43447" heatid="44917" lane="6" entrytime="00:04:15.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.52" />
                    <SPLIT distance="100" swimtime="00:02:11.22" />
                    <SPLIT distance="150" swimtime="00:03:20.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2323" points="177" reactiontime="+122" swimtime="00:01:47.56" resultid="43448" heatid="44926" lane="2" entrytime="00:01:46.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" points="181" reactiontime="+126" swimtime="00:04:06.06" resultid="43449" heatid="45028" lane="5" entrytime="00:04:12.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.52" />
                    <SPLIT distance="100" swimtime="00:02:00.68" />
                    <SPLIT distance="150" swimtime="00:03:06.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernando Manuel" lastname="Pinto" birthdate="1961-05-24" gender="M" nation="POR" license="131365" swrid="5021749" athleteid="43450">
              <RESULTS>
                <RESULT eventid="1058" points="193" swimtime="00:18:01.10" resultid="43451" heatid="45080" lane="1" entrytime="00:17:37.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:02.56" />
                    <SPLIT distance="200" swimtime="00:04:18.47" />
                    <SPLIT distance="300" swimtime="00:06:36.61" />
                    <SPLIT distance="400" swimtime="00:08:55.87" />
                    <SPLIT distance="500" swimtime="00:11:15.68" />
                    <SPLIT distance="600" swimtime="00:13:34.64" />
                    <SPLIT distance="700" swimtime="00:15:50.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2622" points="216" reactiontime="+101" swimtime="00:04:44.35" resultid="43452" heatid="44873" lane="6" entrytime="00:04:44.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.91" />
                    <SPLIT distance="100" swimtime="00:02:18.60" />
                    <SPLIT distance="150" swimtime="00:03:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="192" reactiontime="+108" swimtime="00:08:39.26" resultid="43453" heatid="45124" lane="5" entrytime="00:08:25.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.28" />
                    <SPLIT distance="100" swimtime="00:01:56.64" />
                    <SPLIT distance="150" swimtime="00:03:03.46" />
                    <SPLIT distance="200" swimtime="00:04:11.28" />
                    <SPLIT distance="250" swimtime="00:05:20.91" />
                    <SPLIT distance="300" swimtime="00:06:28.82" />
                    <SPLIT distance="350" swimtime="00:07:36.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Fatima" lastname="Cabral" birthdate="1949-05-20" gender="F" nation="POR" license="106203" swrid="5048947" athleteid="43224">
              <RESULTS>
                <RESULT comment="708 - Não efectuou o ciclo completo de braçada seguida de pernada - SW 7.2" eventid="2173" status="DSQ" swimtime="00:08:03.04" resultid="43225" heatid="45086" lane="6" entrytime="00:07:31.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:01.07" />
                    <SPLIT distance="100" swimtime="00:04:07.50" />
                    <SPLIT distance="150" swimtime="00:06:09.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="65" swimtime="00:01:43.62" resultid="43226" heatid="45097" lane="7" entrytime="00:01:31.28" entrycourse="LCM" />
                <RESULT eventid="2637" points="42" swimtime="00:03:34.83" resultid="43227" heatid="44951" lane="3" entrytime="00:03:18.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:47.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="98" swimtime="00:03:39.29" resultid="43228" heatid="45118" lane="8" entrytime="00:03:29.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:47.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="37" swimtime="00:01:40.14" resultid="43229" heatid="45065" lane="3" entrytime="00:01:26.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cristiano Amaro" lastname="Coelho" birthdate="1988-10-15" gender="M" nation="POR" license="103153" swrid="5231504" athleteid="43268">
              <RESULTS>
                <RESULT eventid="1058" points="329" swimtime="00:11:47.34" resultid="43269" heatid="45084" lane="3" entrytime="00:11:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.37" />
                    <SPLIT distance="200" swimtime="00:02:50.62" />
                    <SPLIT distance="300" swimtime="00:04:20.51" />
                    <SPLIT distance="400" swimtime="00:05:51.15" />
                    <SPLIT distance="500" swimtime="00:07:23.55" />
                    <SPLIT distance="600" swimtime="00:08:55.04" />
                    <SPLIT distance="700" swimtime="00:10:24.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="43270" heatid="45047" lane="3" entrytime="00:00:26.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nuno Manuel" lastname="Sa" birthdate="1971-07-31" gender="M" nation="POR" license="201376" swrid="5171517" athleteid="43501">
              <RESULTS>
                <RESULT eventid="2537" points="288" reactiontime="+88" swimtime="00:01:39.65" resultid="43502" heatid="44885" lane="5" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="315" reactiontime="+87" swimtime="00:03:07.03" resultid="43503" heatid="45093" lane="7" entrytime="00:02:47.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                    <SPLIT distance="100" swimtime="00:01:25.88" />
                    <SPLIT distance="150" swimtime="00:02:16.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="319" reactiontime="+95" swimtime="00:03:36.86" resultid="43504" heatid="44917" lane="5" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.87" />
                    <SPLIT distance="100" swimtime="00:01:47.91" />
                    <SPLIT distance="150" swimtime="00:02:44.11" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="403 - Falsa partida - SW 4.4" eventid="2415" reactiontime="+72" status="DSQ" swimtime="00:01:19.43" resultid="43505" heatid="45109" lane="5" entrytime="00:01:14.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="354" reactiontime="+115" swimtime="00:00:42.06" resultid="43506" heatid="45017" lane="8" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ruben Miguel" lastname="Leodoro" birthdate="1992-10-13" gender="M" nation="POR" license="23484" swrid="4575065" athleteid="43338">
              <RESULTS>
                <RESULT eventid="2537" points="440" reactiontime="+59" swimtime="00:01:17.87" resultid="43339" heatid="44888" lane="5" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="346" reactiontime="+65" swimtime="00:02:56.22" resultid="43340" heatid="44921" lane="2" entrytime="00:02:35.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                    <SPLIT distance="100" swimtime="00:01:25.28" />
                    <SPLIT distance="150" swimtime="00:02:11.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="397" reactiontime="+65" swimtime="00:00:36.42" resultid="43341" heatid="45021" lane="4" entrytime="00:00:33.00" />
                <RESULT eventid="2248" points="362" reactiontime="+83" swimtime="00:06:40.31" resultid="43342" heatid="45061" lane="3" entrytime="00:06:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                    <SPLIT distance="100" swimtime="00:01:29.80" />
                    <SPLIT distance="150" swimtime="00:02:21.12" />
                    <SPLIT distance="200" swimtime="00:03:11.84" />
                    <SPLIT distance="250" swimtime="00:04:11.24" />
                    <SPLIT distance="300" swimtime="00:05:09.75" />
                    <SPLIT distance="350" swimtime="00:05:57.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique Luis" lastname="Seabra" birthdate="1961-04-01" gender="M" nation="POR" license="125467" swrid="4812845" athleteid="43518">
              <RESULTS>
                <RESULT eventid="1058" points="571" swimtime="00:12:33.94" resultid="43519" heatid="45083" lane="7" entrytime="00:12:44.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.90" />
                    <SPLIT distance="300" swimtime="00:04:30.64" />
                    <SPLIT distance="400" swimtime="00:06:06.80" />
                    <SPLIT distance="500" swimtime="00:07:42.54" />
                    <SPLIT distance="600" swimtime="00:09:19.98" />
                    <SPLIT distance="700" swimtime="00:10:57.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="554" reactiontime="+82" swimtime="00:02:50.31" resultid="43520" heatid="45093" lane="2" entrytime="00:02:47.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                    <SPLIT distance="100" swimtime="00:01:16.29" />
                    <SPLIT distance="150" swimtime="00:02:02.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="433" reactiontime="+87" swimtime="00:03:30.15" resultid="43521" heatid="44977" lane="7" entrytime="00:03:32.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                    <SPLIT distance="100" swimtime="00:01:41.92" />
                    <SPLIT distance="150" swimtime="00:02:43.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="511" reactiontime="+85" swimtime="00:06:14.89" resultid="43522" heatid="45128" lane="3" entrytime="00:06:07.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:19.50" />
                    <SPLIT distance="150" swimtime="00:02:03.63" />
                    <SPLIT distance="200" swimtime="00:02:50.55" />
                    <SPLIT distance="250" swimtime="00:03:38.83" />
                    <SPLIT distance="300" swimtime="00:04:29.79" />
                    <SPLIT distance="350" swimtime="00:05:21.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="444" reactiontime="+103" swimtime="00:07:33.45" resultid="43523" heatid="45059" lane="5" entrytime="00:07:47.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.54" />
                    <SPLIT distance="100" swimtime="00:01:45.90" />
                    <SPLIT distance="150" swimtime="00:02:55.50" />
                    <SPLIT distance="200" swimtime="00:04:05.37" />
                    <SPLIT distance="250" swimtime="00:05:03.97" />
                    <SPLIT distance="300" swimtime="00:06:03.62" />
                    <SPLIT distance="350" swimtime="00:06:48.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ines Silva" lastname="Carvalho" birthdate="1983-08-16" gender="F" nation="POR" license="212606" swrid="5429040" athleteid="43244">
              <RESULTS>
                <RESULT eventid="1060" points="184" swimtime="00:17:01.67" resultid="43245" heatid="45075" lane="8" entrytime="00:18:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:04:09.35" />
                    <SPLIT distance="200" swimtime="00:06:19.60" />
                    <SPLIT distance="400" swimtime="00:08:29.63" />
                    <SPLIT distance="500" swimtime="00:10:37.48" />
                    <SPLIT distance="600" swimtime="00:12:47.88" />
                    <SPLIT distance="700" swimtime="00:14:59.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2173" points="324" swimtime="00:03:51.37" resultid="43246" heatid="45088" lane="2" entrytime="00:03:55.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.03" />
                    <SPLIT distance="100" swimtime="00:01:53.71" />
                    <SPLIT distance="150" swimtime="00:02:53.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="285" reactiontime="+96" swimtime="00:01:50.25" resultid="43247" heatid="45121" lane="1" entrytime="00:01:47.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="178" reactiontime="+102" swimtime="00:08:18.80" resultid="43248" heatid="45008" lane="3" entrytime="00:09:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.45" />
                    <SPLIT distance="100" swimtime="00:01:58.52" />
                    <SPLIT distance="150" swimtime="00:03:00.96" />
                    <SPLIT distance="200" swimtime="00:04:04.82" />
                    <SPLIT distance="250" swimtime="00:05:08.09" />
                    <SPLIT distance="300" swimtime="00:06:12.96" />
                    <SPLIT distance="350" swimtime="00:07:16.03" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="809 - Movimento alternado de pernas durante o percurso - SW 8.3" eventid="2667" reactiontime="+106" status="DSQ" swimtime="00:04:23.76" resultid="43249" heatid="45031" lane="2" entrytime="00:04:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.34" />
                    <SPLIT distance="100" swimtime="00:02:04.62" />
                    <SPLIT distance="150" swimtime="00:03:13.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Pedro" lastname="Neves" birthdate="1981-09-08" gender="M" nation="POR" license="17203" swrid="4190112" athleteid="43402">
              <RESULTS>
                <RESULT eventid="2415" status="DNS" swimtime="00:00:00.00" resultid="43403" heatid="45115" lane="7" entrytime="00:01:00.17" entrycourse="SCM" />
                <RESULT eventid="2263" status="DNS" swimtime="00:00:00.00" resultid="43404" heatid="45131" lane="3" entrytime="00:04:45.82" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena Maria" lastname="Cardoso" birthdate="1966-08-26" gender="F" nation="POR" license="205207" swrid="5231500" athleteid="43233">
              <RESULTS>
                <RESULT eventid="1060" points="164" swimtime="00:18:25.03" resultid="43234" heatid="45075" lane="1" entrytime="00:17:35.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:02.94" />
                    <SPLIT distance="200" swimtime="00:04:20.92" />
                    <SPLIT distance="300" swimtime="00:06:43.25" />
                    <SPLIT distance="400" swimtime="00:09:04.70" />
                    <SPLIT distance="500" swimtime="00:11:24.97" />
                    <SPLIT distance="600" swimtime="00:13:45.46" />
                    <SPLIT distance="700" swimtime="00:16:07.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2203" points="259" reactiontime="+132" swimtime="00:02:02.51" resultid="43235" heatid="44881" lane="8" entrytime="00:02:01.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2308" points="254" reactiontime="+136" swimtime="00:04:23.51" resultid="43236" heatid="44913" lane="7" entrytime="00:04:26.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.60" />
                    <SPLIT distance="100" swimtime="00:02:04.71" />
                    <SPLIT distance="150" swimtime="00:03:14.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="250" reactiontime="+156" swimtime="00:00:56.68" resultid="43237" heatid="45023" lane="3" entrytime="00:01:01.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jaime Alberto" lastname="Milheiro" birthdate="1970-12-20" gender="M" nation="POR" license="16023" swrid="4558725" athleteid="43381">
              <RESULTS>
                <RESULT eventid="2682" points="591" reactiontime="+94" swimtime="00:00:32.92" resultid="43382" heatid="44898" lane="2" entrytime="00:00:31.59" entrycourse="SCM" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="43383" heatid="45044" lane="6" entrytime="00:00:28.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabel Maria" lastname="Pinto" birthdate="1972-02-03" gender="F" nation="POR" license="207697" swrid="5292300" athleteid="43454">
              <RESULTS>
                <RESULT eventid="1060" points="196" swimtime="00:16:38.91" resultid="43455" heatid="45074" lane="2" entrytime="00:19:20.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:57.06" />
                    <SPLIT distance="200" swimtime="00:04:01.92" />
                    <SPLIT distance="300" swimtime="00:06:08.54" />
                    <SPLIT distance="400" swimtime="00:08:15.81" />
                    <SPLIT distance="500" swimtime="00:10:22.82" />
                    <SPLIT distance="600" swimtime="00:12:29.83" />
                    <SPLIT distance="700" swimtime="00:14:37.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2203" points="176" reactiontime="+119" swimtime="00:02:05.56" resultid="43456" heatid="44880" lane="5" entrytime="00:02:02.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2308" points="215" reactiontime="+122" swimtime="00:04:25.46" resultid="43457" heatid="44913" lane="6" entrytime="00:04:15.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.30" />
                    <SPLIT distance="100" swimtime="00:02:11.86" />
                    <SPLIT distance="150" swimtime="00:03:23.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="189" reactiontime="+105" swimtime="00:00:54.59" resultid="43458" heatid="45024" lane="2" entrytime="00:00:53.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo Sergio" lastname="Pereira" birthdate="1974-04-20" gender="M" nation="POR" license="153326" swrid="5117187" athleteid="43440">
              <RESULTS>
                <RESULT eventid="2622" status="DNS" swimtime="00:00:00.00" resultid="43441" heatid="44877" lane="7" entrytime="00:03:20.00" />
                <RESULT eventid="2188" status="DNS" swimtime="00:00:00.00" resultid="43442" heatid="44945" lane="4" entrytime="00:00:41.91" entrycourse="LCM" />
                <RESULT eventid="2445" status="DNS" swimtime="00:00:00.00" resultid="43443" heatid="44996" lane="4" entrytime="00:01:30.20" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Manuel" lastname="Pinto" birthdate="1979-01-21" gender="M" nation="POR" license="106876" swrid="4598766" athleteid="43459">
              <RESULTS>
                <RESULT eventid="2218" points="400" reactiontime="+96" swimtime="00:03:01.57" resultid="43460" heatid="44920" lane="5" entrytime="00:02:52.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                    <SPLIT distance="100" swimtime="00:01:27.94" />
                    <SPLIT distance="150" swimtime="00:02:16.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2323" points="300" reactiontime="+94" swimtime="00:01:27.61" resultid="43461" heatid="44927" lane="7" entrytime="00:01:22.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="428" reactiontime="+89" swimtime="00:01:12.04" resultid="43462" heatid="45108" lane="3" entrytime="00:01:18.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="305" reactiontime="+106" swimtime="00:03:16.68" resultid="43463" heatid="44980" lane="4" entrytime="00:02:49.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                    <SPLIT distance="100" swimtime="00:01:28.63" />
                    <SPLIT distance="150" swimtime="00:02:26.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" status="DNS" swimtime="00:00:00.00" resultid="43464" heatid="45030" lane="8" entrytime="00:03:11.58" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nuno Silva" lastname="Lobo" birthdate="1963-12-13" gender="M" nation="POR" license="102544" swrid="5036815" athleteid="43343">
              <RESULTS>
                <RESULT eventid="2567" points="322" reactiontime="+111" swimtime="00:03:46.19" resultid="43344" heatid="45029" lane="7" entrytime="00:03:42.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.51" />
                    <SPLIT distance="100" swimtime="00:01:48.28" />
                    <SPLIT distance="150" swimtime="00:02:47.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="612" reactiontime="+80" swimtime="00:02:57.75" resultid="43345" heatid="44919" lane="3" entrytime="00:03:15.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                    <SPLIT distance="100" swimtime="00:01:27.82" />
                    <SPLIT distance="150" swimtime="00:02:12.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="670" reactiontime="+90" swimtime="00:02:55.03" resultid="43346" heatid="44978" lane="4" entrytime="00:03:09.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="100" swimtime="00:01:22.35" />
                    <SPLIT distance="150" swimtime="00:02:14.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="642" reactiontime="+72" swimtime="00:00:36.29" resultid="43347" heatid="45019" lane="4" entrytime="00:00:36.95" entrycourse="LCM" />
                <RESULT eventid="2248" points="580" reactiontime="+111" swimtime="00:06:36.95" resultid="43348" heatid="45061" lane="8" entrytime="00:06:31.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                    <SPLIT distance="100" swimtime="00:01:40.25" />
                    <SPLIT distance="150" swimtime="00:02:34.91" />
                    <SPLIT distance="200" swimtime="00:03:26.13" />
                    <SPLIT distance="250" swimtime="00:04:20.79" />
                    <SPLIT distance="300" swimtime="00:05:16.17" />
                    <SPLIT distance="350" swimtime="00:05:58.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabel Carolina" lastname="Neves" birthdate="1980-03-27" gender="F" nation="POR" license="202850" swrid="4889296" athleteid="43396">
              <RESULTS>
                <RESULT eventid="1060" points="312" swimtime="00:14:26.23" resultid="43397" heatid="45076" lane="3" entrytime="00:14:33.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.61" />
                    <SPLIT distance="200" swimtime="00:03:26.70" />
                    <SPLIT distance="300" swimtime="00:05:16.71" />
                    <SPLIT distance="400" swimtime="00:07:07.99" />
                    <SPLIT distance="500" swimtime="00:09:00.82" />
                    <SPLIT distance="600" swimtime="00:10:53.24" />
                    <SPLIT distance="700" swimtime="00:12:42.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2278" points="314" reactiontime="+106" swimtime="00:03:13.61" resultid="43398" heatid="44903" lane="5" entrytime="00:03:10.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.29" />
                    <SPLIT distance="100" swimtime="00:01:32.86" />
                    <SPLIT distance="150" swimtime="00:02:25.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2308" points="243" reactiontime="+88" swimtime="00:04:06.43" resultid="43399" heatid="44914" lane="7" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.65" />
                    <SPLIT distance="100" swimtime="00:02:04.24" />
                    <SPLIT distance="150" swimtime="00:03:07.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="304" reactiontime="+95" swimtime="00:07:00.35" resultid="43400" heatid="45010" lane="5" entrytime="00:07:08.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.18" />
                    <SPLIT distance="100" swimtime="00:01:37.35" />
                    <SPLIT distance="150" swimtime="00:02:32.23" />
                    <SPLIT distance="200" swimtime="00:03:26.31" />
                    <SPLIT distance="250" swimtime="00:04:21.63" />
                    <SPLIT distance="300" swimtime="00:05:15.50" />
                    <SPLIT distance="350" swimtime="00:06:08.52" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="604 - Durante o percurso perdeu a posição dorsal - SW 6.2" eventid="2400" reactiontime="+111" status="DSQ" swimtime="00:08:58.82" resultid="43401" heatid="45064" lane="1" entrytime="00:08:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.34" />
                    <SPLIT distance="100" swimtime="00:01:59.50" />
                    <SPLIT distance="150" swimtime="00:03:27.43" />
                    <SPLIT distance="200" swimtime="00:04:30.40" />
                    <SPLIT distance="250" swimtime="00:05:49.24" />
                    <SPLIT distance="300" swimtime="00:07:06.47" />
                    <SPLIT distance="350" swimtime="00:08:04.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Teresa" lastname="Brandao" birthdate="1969-05-11" gender="F" nation="POR" license="108037" swrid="4319543" athleteid="43218">
              <RESULTS>
                <RESULT eventid="2552" points="497" reactiontime="+99" swimtime="00:01:30.19" resultid="43219" heatid="44924" lane="1" entrytime="00:01:28.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="555" swimtime="00:12:00.70" resultid="43220" heatid="45078" lane="6" entrytime="00:11:41.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.82" />
                    <SPLIT distance="200" swimtime="00:02:49.64" />
                    <SPLIT distance="300" swimtime="00:04:19.82" />
                    <SPLIT distance="400" swimtime="00:05:52.06" />
                    <SPLIT distance="500" swimtime="00:07:25.47" />
                    <SPLIT distance="600" swimtime="00:08:57.94" />
                    <SPLIT distance="700" swimtime="00:10:30.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2278" points="648" reactiontime="+96" swimtime="00:02:39.50" resultid="43221" heatid="44905" lane="1" entrytime="00:02:38.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                    <SPLIT distance="100" swimtime="00:01:17.35" />
                    <SPLIT distance="150" swimtime="00:01:58.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="552" reactiontime="+108" swimtime="00:05:51.43" resultid="43222" heatid="45013" lane="1" entrytime="00:05:44.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                    <SPLIT distance="100" swimtime="00:01:24.32" />
                    <SPLIT distance="150" swimtime="00:02:08.16" />
                    <SPLIT distance="200" swimtime="00:02:53.43" />
                    <SPLIT distance="250" swimtime="00:03:38.29" />
                    <SPLIT distance="300" swimtime="00:04:23.15" />
                    <SPLIT distance="350" swimtime="00:05:08.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2400" points="485" reactiontime="+101" swimtime="00:07:04.98" resultid="43223" heatid="45064" lane="6" entrytime="00:06:46.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.97" />
                    <SPLIT distance="100" swimtime="00:01:39.98" />
                    <SPLIT distance="150" swimtime="00:02:36.90" />
                    <SPLIT distance="200" swimtime="00:03:32.96" />
                    <SPLIT distance="250" swimtime="00:04:34.37" />
                    <SPLIT distance="300" swimtime="00:05:34.88" />
                    <SPLIT distance="350" swimtime="00:06:21.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Catarina Bayer" lastname="Castro" birthdate="1973-10-11" gender="F" nation="POR" license="127874" swrid="4905768" athleteid="43250">
              <RESULTS>
                <RESULT eventid="2552" points="277" reactiontime="+111" swimtime="00:01:43.89" resultid="43251" heatid="44923" lane="3" entrytime="00:01:46.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="319" reactiontime="+110" swimtime="00:03:42.41" resultid="43252" heatid="44972" lane="1" entrytime="00:03:47.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.94" />
                    <SPLIT distance="100" swimtime="00:01:48.12" />
                    <SPLIT distance="150" swimtime="00:02:53.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="247" reactiontime="+128" swimtime="00:00:49.95" resultid="43253" heatid="45023" lane="4" entrytime="00:00:57.77" entrycourse="LCM" />
                <RESULT eventid="2667" points="319" reactiontime="+112" swimtime="00:03:47.71" resultid="43254" heatid="45031" lane="6" entrytime="00:03:57.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.96" />
                    <SPLIT distance="100" swimtime="00:01:47.93" />
                    <SPLIT distance="150" swimtime="00:02:47.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2400" points="344" reactiontime="+107" swimtime="00:07:54.62" resultid="43255" heatid="45064" lane="8" entrytime="00:08:18.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.68" />
                    <SPLIT distance="100" swimtime="00:01:49.32" />
                    <SPLIT distance="150" swimtime="00:02:51.08" />
                    <SPLIT distance="200" swimtime="00:03:53.42" />
                    <SPLIT distance="250" swimtime="00:05:04.80" />
                    <SPLIT distance="300" swimtime="00:06:13.20" />
                    <SPLIT distance="350" swimtime="00:07:03.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel Pinheiro" lastname="Pires" birthdate="1978-08-05" gender="M" nation="POR" license="153288" swrid="5115795" athleteid="43465">
              <RESULTS>
                <RESULT eventid="2323" points="638" reactiontime="+69" swimtime="00:01:08.14" resultid="43466" heatid="44930" lane="2" entrytime="00:01:04.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="684" reactiontime="+73" swimtime="00:01:01.65" resultid="43467" heatid="45104" lane="6" entrytime="00:01:00.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" status="DNS" swimtime="00:00:00.00" resultid="43468" heatid="44981" lane="2" entrytime="00:02:45.00" />
                <RESULT eventid="2293" points="554" reactiontime="+62" swimtime="00:00:34.56" resultid="43469" heatid="45021" lane="2" entrytime="00:00:33.00" />
                <RESULT eventid="2652" points="707" reactiontime="+63" swimtime="00:00:27.58" resultid="43470" heatid="45047" lane="8" entrytime="00:00:27.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo Francisco" lastname="Torres" birthdate="1962-11-12" gender="M" nation="POR" license="130665" swrid="5001750" athleteid="43554">
              <RESULTS>
                <RESULT eventid="2263" status="DNS" swimtime="00:00:00.00" resultid="43555" heatid="45129" lane="5" entrytime="00:05:42.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Regina" lastname="Mendes" birthdate="1965-01-01" gender="F" nation="POR" license="26842" swrid="4575257" athleteid="43372">
              <RESULTS>
                <RESULT eventid="2233" status="DNS" swimtime="00:00:00.00" resultid="43373" heatid="44972" lane="2" entrytime="00:03:37.49" entrycourse="LCM" />
                <RESULT eventid="2460" status="DNS" swimtime="00:00:00.00" resultid="43374" heatid="45121" lane="2" entrytime="00:01:45.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Maria" lastname="Cunha" birthdate="1971-09-03" gender="M" nation="POR" license="204079" swrid="4548183" athleteid="43285">
              <RESULTS>
                <RESULT eventid="2652" points="436" reactiontime="+124" swimtime="00:00:33.11" resultid="43286" heatid="45039" lane="7" entrytime="00:00:33.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Augusto" lastname="Vaz" birthdate="1965-09-27" gender="M" nation="POR" license="133405" swrid="5090073" athleteid="43562">
              <RESULTS>
                <RESULT eventid="2682" points="693" reactiontime="+73" swimtime="00:00:31.96" resultid="43563" heatid="44898" lane="8" entrytime="00:00:32.59" entrycourse="LCM" />
                <RESULT eventid="2188" points="632" reactiontime="+77" swimtime="00:00:36.18" resultid="43564" heatid="44949" lane="2" entrytime="00:00:35.55" entrycourse="LCM" />
                <RESULT comment="Rec Nac Esc G" eventid="2445" points="707" reactiontime="+76" swimtime="00:01:21.51" resultid="43565" heatid="44998" lane="5" entrytime="00:01:19.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="532" reactiontime="+75" swimtime="00:00:38.63" resultid="43566" heatid="45019" lane="7" entrytime="00:00:39.29" entrycourse="LCM" />
                <RESULT comment="403 - Falsa partida - SW 4.4" eventid="2652" reactiontime="+65" status="DSQ" swimtime="00:00:29.57" resultid="43567" heatid="45044" lane="2" entrytime="00:00:28.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo Jorge" lastname="Rocha" birthdate="1959-05-22" gender="M" nation="POR" license="208405" swrid="5326942" athleteid="43487">
              <RESULTS>
                <RESULT eventid="1058" points="309" swimtime="00:15:25.19" resultid="43488" heatid="45081" lane="7" entrytime="00:15:31.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.38" />
                    <SPLIT distance="200" swimtime="00:03:46.59" />
                    <SPLIT distance="300" swimtime="00:05:44.32" />
                    <SPLIT distance="400" swimtime="00:07:43.39" />
                    <SPLIT distance="500" swimtime="00:09:41.28" />
                    <SPLIT distance="600" swimtime="00:11:39.19" />
                    <SPLIT distance="700" swimtime="00:13:36.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2622" points="265" reactiontime="+148" swimtime="00:04:25.59" resultid="43489" heatid="44874" lane="6" entrytime="00:04:03.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.71" />
                    <SPLIT distance="100" swimtime="00:02:09.45" />
                    <SPLIT distance="150" swimtime="00:03:22.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="295" reactiontime="+134" swimtime="00:03:29.96" resultid="43490" heatid="45091" lane="8" entrytime="00:03:38.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.94" />
                    <SPLIT distance="100" swimtime="00:01:40.03" />
                    <SPLIT distance="150" swimtime="00:02:36.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="308" reactiontime="+142" swimtime="00:07:23.81" resultid="43491" heatid="45126" lane="1" entrytime="00:07:34.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.11" />
                    <SPLIT distance="100" swimtime="00:01:40.82" />
                    <SPLIT distance="150" swimtime="00:02:37.54" />
                    <SPLIT distance="200" swimtime="00:03:36.31" />
                    <SPLIT distance="250" swimtime="00:04:33.43" />
                    <SPLIT distance="300" swimtime="00:05:33.08" />
                    <SPLIT distance="350" swimtime="00:06:32.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CNMAIA" nation="POR" region="ANNP" clubid="42667" swrid="65883" name="Clube de Natacao da Maia" shortname="Natacao da Maia">
          <ATHLETES>
            <ATHLETE firstname="Jose Luis" lastname="Moreira" birthdate="1993-07-22" gender="M" nation="POR" license="207903" swrid="5065717" athleteid="42682">
              <RESULTS>
                <RESULT eventid="2622" points="436" reactiontime="+83" swimtime="00:03:10.78" resultid="42683" heatid="44877" lane="3" entrytime="00:03:18.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                    <SPLIT distance="100" swimtime="00:01:30.83" />
                    <SPLIT distance="150" swimtime="00:02:20.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="354" reactiontime="+90" swimtime="00:00:35.43" resultid="42684" heatid="44896" lane="7" entrytime="00:00:36.79" entrycourse="LCM" />
                <RESULT eventid="2188" points="472" reactiontime="+80" swimtime="00:00:37.07" resultid="42685" heatid="44946" lane="5" entrytime="00:00:39.92" entrycourse="LCM" />
                <RESULT eventid="2415" points="462" reactiontime="+80" swimtime="00:01:06.87" resultid="42686" heatid="45110" lane="5" entrytime="00:01:10.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="489" reactiontime="+77" swimtime="00:00:29.38" resultid="42687" heatid="45043" lane="7" entrytime="00:00:29.22" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Pedro" lastname="Ferreira" birthdate="1995-12-25" gender="M" nation="POR" license="111411" swrid="4398286" athleteid="42673">
              <RESULTS>
                <RESULT eventid="2537" points="427" reactiontime="+59" swimtime="00:01:18.67" resultid="42674" heatid="44886" lane="2" entrytime="00:01:34.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="458" reactiontime="+78" swimtime="00:00:32.52" resultid="42675" heatid="44897" lane="3" entrytime="00:00:33.33" />
                <RESULT eventid="2323" points="389" reactiontime="+78" swimtime="00:01:17.84" resultid="42676" heatid="44928" lane="1" entrytime="00:01:13.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="381" reactiontime="+80" swimtime="00:02:53.77" resultid="42677" heatid="44979" lane="6" entrytime="00:02:58.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="100" swimtime="00:01:20.73" />
                    <SPLIT distance="150" swimtime="00:02:13.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="403" reactiontime="+60" swimtime="00:00:36.24" resultid="42678" heatid="45019" lane="2" entrytime="00:00:39.15" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Goncalves" lastname="Oliveira" birthdate="1993-09-07" gender="M" nation="POR" license="20359" swrid="4575419" athleteid="42699">
              <RESULTS>
                <RESULT eventid="2537" points="738" reactiontime="+61" swimtime="00:01:05.56" resultid="42700" heatid="44888" lane="4" entrytime="00:01:04.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="713" reactiontime="+68" swimtime="00:00:28.06" resultid="42701" heatid="44901" lane="6" entrytime="00:00:27.64" entrycourse="LCM" />
                <RESULT eventid="2323" points="750" reactiontime="+73" swimtime="00:01:02.57" resultid="42702" heatid="44930" lane="6" entrytime="00:01:02.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="723" reactiontime="+68" swimtime="00:00:57.59" resultid="42703" heatid="45116" lane="8" entrytime="00:00:57.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="704" reactiontime="+57" swimtime="00:00:30.09" resultid="42704" heatid="45022" lane="4" entrytime="00:00:29.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Manuela" lastname="Neto" birthdate="1962-07-04" gender="F" nation="POR" license="102090" swrid="4319547" athleteid="42688">
              <RESULTS>
                <RESULT eventid="1060" points="252" swimtime="00:15:56.51" resultid="42689" heatid="45075" lane="3" entrytime="00:15:57.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:52.24" />
                    <SPLIT distance="200" swimtime="00:03:54.14" />
                    <SPLIT distance="300" swimtime="00:05:54.15" />
                    <SPLIT distance="400" swimtime="00:07:54.75" />
                    <SPLIT distance="500" swimtime="00:09:55.54" />
                    <SPLIT distance="600" swimtime="00:11:56.26" />
                    <SPLIT distance="700" swimtime="00:13:57.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2278" points="256" swimtime="00:03:40.14" resultid="42690" heatid="44902" lane="6" entrytime="00:03:50.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.95" />
                    <SPLIT distance="100" swimtime="00:01:45.20" />
                    <SPLIT distance="150" swimtime="00:02:43.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="253" swimtime="00:01:40.62" resultid="42691" heatid="44953" lane="3" entrytime="00:01:40.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="264" swimtime="00:07:32.97" resultid="42692" heatid="45009" lane="3" entrytime="00:07:49.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.55" />
                    <SPLIT distance="100" swimtime="00:01:45.71" />
                    <SPLIT distance="150" swimtime="00:02:42.03" />
                    <SPLIT distance="200" swimtime="00:03:42.53" />
                    <SPLIT distance="250" swimtime="00:04:39.33" />
                    <SPLIT distance="300" swimtime="00:05:38.96" />
                    <SPLIT distance="350" swimtime="00:06:36.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="289" swimtime="00:00:44.74" resultid="42693" heatid="45068" lane="8" entrytime="00:00:42.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Manuel" lastname="Ribeiro" birthdate="1969-11-03" gender="M" nation="POR" license="201429" swrid="5171513" athleteid="42705">
              <RESULTS>
                <RESULT eventid="1058" points="263" swimtime="00:14:19.81" resultid="42706" heatid="45082" lane="2" entrytime="00:13:41.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.66" />
                    <SPLIT distance="200" swimtime="00:03:27.30" />
                    <SPLIT distance="300" swimtime="00:05:16.49" />
                    <SPLIT distance="400" swimtime="00:07:06.69" />
                    <SPLIT distance="500" swimtime="00:08:56.82" />
                    <SPLIT distance="600" swimtime="00:10:45.65" />
                    <SPLIT distance="700" swimtime="00:12:33.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Mafalda" lastname="Oliveira" birthdate="1981-03-30" gender="F" nation="POR" license="23193" swrid="4061391" athleteid="42694">
              <RESULTS>
                <RESULT eventid="1060" points="488" swimtime="00:12:26.77" resultid="42695" heatid="45078" lane="8" entrytime="00:12:20.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.98" />
                    <SPLIT distance="200" swimtime="00:02:56.57" />
                    <SPLIT distance="300" swimtime="00:04:31.75" />
                    <SPLIT distance="400" swimtime="00:06:07.37" />
                    <SPLIT distance="500" swimtime="00:07:43.41" />
                    <SPLIT distance="600" swimtime="00:09:17.84" />
                    <SPLIT distance="700" swimtime="00:10:53.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2278" points="458" reactiontime="+80" swimtime="00:02:50.70" resultid="42696" heatid="44905" lane="8" entrytime="00:02:48.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                    <SPLIT distance="100" swimtime="00:01:19.83" />
                    <SPLIT distance="150" swimtime="00:02:05.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="549" reactiontime="+84" swimtime="00:03:04.95" resultid="42697" heatid="44973" lane="5" entrytime="00:03:07.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                    <SPLIT distance="100" swimtime="00:01:25.42" />
                    <SPLIT distance="150" swimtime="00:02:22.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="480" reactiontime="+84" swimtime="00:06:00.99" resultid="42698" heatid="45012" lane="4" entrytime="00:06:05.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.60" />
                    <SPLIT distance="100" swimtime="00:01:23.68" />
                    <SPLIT distance="150" swimtime="00:02:09.26" />
                    <SPLIT distance="200" swimtime="00:02:55.72" />
                    <SPLIT distance="250" swimtime="00:03:42.14" />
                    <SPLIT distance="300" swimtime="00:04:28.56" />
                    <SPLIT distance="350" swimtime="00:05:14.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Pedro" lastname="Ferreira" birthdate="1964-06-30" gender="M" nation="POR" license="129087" swrid="4951641" athleteid="42679">
              <RESULTS>
                <RESULT eventid="2293" points="181" reactiontime="+100" swimtime="00:00:55.27" resultid="42680" heatid="45015" lane="3" entrytime="00:00:56.13" entrycourse="LCM" />
                <RESULT eventid="2652" points="332" reactiontime="+99" swimtime="00:00:38.41" resultid="42681" heatid="45036" lane="7" entrytime="00:00:37.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Pedro" lastname="Bandeira" birthdate="1995-12-20" gender="M" nation="POR" license="24291" swrid="4123339" athleteid="42668">
              <RESULTS>
                <RESULT eventid="2188" points="621" reactiontime="+71" swimtime="00:00:33.85" resultid="42669" heatid="44947" lane="7" entrytime="00:00:39.28" />
                <RESULT eventid="2652" points="575" reactiontime="+64" swimtime="00:00:27.84" resultid="42670" heatid="45041" lane="6" entrytime="00:00:31.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo Jorge" lastname="Corado" birthdate="1967-05-30" gender="M" nation="POR" license="206893" swrid="5276310" athleteid="42671">
              <RESULTS>
                <RESULT eventid="2652" points="215" reactiontime="+124" swimtime="00:00:41.87" resultid="42672" heatid="45033" lane="4" entrytime="00:00:46.56" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ADRCIMM" nation="POR" region="ANL" clubid="41793" swrid="86260" name="Assoc Desp Rec Colegio Int Monte Maior" shortname="Colegio Monte Maior">
          <ATHLETES>
            <ATHLETE firstname="Jorge Miguel" lastname="Silva" birthdate="1976-01-15" gender="M" nation="POR" license="119954" swrid="4614048" athleteid="41794">
              <RESULTS>
                <RESULT eventid="2415" status="DNS" swimtime="00:00:00.00" resultid="41795" heatid="45110" lane="4" entrytime="00:01:10.00" />
                <RESULT eventid="2445" status="DNS" swimtime="00:00:00.00" resultid="41796" heatid="44997" lane="8" entrytime="00:01:30.00" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CNLX" nation="POR" region="ANL" clubid="42321" swrid="90828" name="Clube de Natacao de Lisboa" shortname="Natacao de Lisboa">
          <ATHLETES>
            <ATHLETE firstname="Laura" lastname="Pola" birthdate="1992-05-06" gender="F" nation="ITA" license="214291" athleteid="42349">
              <RESULTS>
                <RESULT eventid="2338" status="DNS" swimtime="00:00:00.00" resultid="42350" heatid="44890" lane="3" entrytime="00:00:45.00" />
                <RESULT eventid="2278" points="474" reactiontime="+86" swimtime="00:02:43.75" resultid="42351" heatid="44903" lane="6" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:16.14" />
                    <SPLIT distance="150" swimtime="00:01:59.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="510" reactiontime="+95" swimtime="00:01:11.63" resultid="42352" heatid="44954" lane="5" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="527" reactiontime="+84" swimtime="00:00:32.31" resultid="42353" heatid="45070" lane="7" entrytime="00:00:36.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rodrigo Serra" lastname="Farias" birthdate="1996-10-29" gender="M" nation="POR" license="106392" swrid="4285282" athleteid="42322">
              <RESULTS>
                <RESULT eventid="2682" points="789" reactiontime="+69" swimtime="00:00:27.13" resultid="42323" heatid="44901" lane="5" entrytime="00:00:27.00" />
                <RESULT eventid="2507" points="629" reactiontime="+68" swimtime="00:02:14.37" resultid="42324" heatid="45096" lane="3" entrytime="00:02:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                    <SPLIT distance="100" swimtime="00:01:05.41" />
                    <SPLIT distance="150" swimtime="00:01:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2323" points="727" reactiontime="+72" swimtime="00:01:03.23" resultid="42325" heatid="44930" lane="3" entrytime="00:01:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="745" reactiontime="+68" swimtime="00:00:57.04" resultid="42326" heatid="45116" lane="5" entrytime="00:00:55.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" status="WDR" swimtime="00:00:00.00" resultid="42327" entrytime="00:02:25.00" />
                <RESULT eventid="2652" points="735" reactiontime="+68" swimtime="00:00:25.65" resultid="42328" heatid="45048" lane="4" entrytime="00:00:25.02" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno Calado" lastname="Camara" birthdate="1977-04-18" gender="M" nation="POR" license="128759" swrid="4934088" athleteid="42335">
              <RESULTS>
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="42336" heatid="45046" lane="3" entrytime="00:00:27.43" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre Filipe" lastname="Carocha" birthdate="1994-08-26" gender="M" nation="POR" license="127747" swrid="4905792" athleteid="42337">
              <RESULTS>
                <RESULT eventid="2682" status="DNS" swimtime="00:00:00.00" resultid="42338" heatid="44901" lane="1" entrytime="00:00:28.40" />
                <RESULT eventid="2507" status="WDR" swimtime="00:00:00.00" resultid="42339" entrytime="00:02:15.00" />
                <RESULT eventid="2323" status="DNS" swimtime="00:00:00.00" resultid="42340" heatid="44929" lane="4" entrytime="00:01:05.29" />
                <RESULT eventid="2415" status="DNS" swimtime="00:00:00.00" resultid="42341" heatid="45116" lane="3" entrytime="00:00:55.78" />
                <RESULT eventid="2293" status="DNS" swimtime="00:00:00.00" resultid="42342" heatid="45022" lane="8" entrytime="00:00:32.98" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="42343" heatid="45048" lane="6" entrytime="00:00:25.68" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rita Fernandes" lastname="Leitao" birthdate="1996-08-29" gender="F" nation="POR" license="25571" swrid="4561991" athleteid="42329">
              <RESULTS>
                <RESULT eventid="2173" points="703" swimtime="00:02:55.23" resultid="42330" heatid="45089" lane="4" entrytime="00:02:40.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:01:22.72" />
                    <SPLIT distance="150" swimtime="00:02:08.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="741" reactiontime="+82" swimtime="00:00:36.07" resultid="42331" heatid="45103" lane="5" entrytime="00:00:36.19" />
                <RESULT comment="Rec Nac Esc A" eventid="2637" points="759" reactiontime="+80" swimtime="00:01:02.77" resultid="42332" heatid="44957" lane="4" entrytime="00:01:00.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="806" reactiontime="+80" swimtime="00:01:17.74" resultid="42333" heatid="45123" lane="5" entrytime="00:01:19.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="731" reactiontime="+76" swimtime="00:00:28.97" resultid="42334" heatid="45073" lane="4" entrytime="00:00:28.77" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Claudia Alexandra" lastname="Mendes" birthdate="1995-05-05" gender="F" nation="POR" license="126614" swrid="4860214" athleteid="42344">
              <RESULTS>
                <RESULT eventid="2522" points="489" reactiontime="+69" swimtime="00:00:38.78" resultid="42345" heatid="45027" lane="6" entrytime="00:00:36.15" />
                <RESULT eventid="2430" points="472" reactiontime="+94" swimtime="00:00:33.51" resultid="42346" heatid="45072" lane="2" entrytime="00:00:31.57" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Maria" lastname="Rosa" birthdate="1991-11-15" gender="M" nation="POR" license="25532" swrid="4559955" athleteid="42347">
              <RESULTS>
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="42348" heatid="45042" lane="4" entrytime="00:00:29.50" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="PORTIN" nation="POR" region="ANALG" clubid="42707" swrid="65802" name="Portinado-Assoc Natacao de Portimao" shortname="Portinado">
          <ATHLETES>
            <ATHLETE firstname="Adriana Pereira" lastname="Valentim" birthdate="1992-04-15" gender="F" nation="POR" license="13347" swrid="4074228" athleteid="42735">
              <RESULTS>
                <RESULT eventid="2203" points="596" reactiontime="+81" swimtime="00:01:19.00" resultid="42736" heatid="44883" lane="3" entrytime="00:01:17.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2338" points="508" reactiontime="+94" swimtime="00:00:34.82" resultid="42737" heatid="44891" lane="3" entrytime="00:00:36.84" />
                <RESULT eventid="2607" points="525" reactiontime="+86" swimtime="00:00:40.47" resultid="42738" heatid="45103" lane="1" entrytime="00:00:41.62" entrycourse="LCM" />
                <RESULT eventid="2522" points="651" reactiontime="+70" swimtime="00:00:35.26" resultid="42739" heatid="45027" lane="3" entrytime="00:00:34.13" entrycourse="LCM" />
                <RESULT eventid="2430" points="602" reactiontime="+83" swimtime="00:00:30.90" resultid="42740" heatid="45071" lane="3" entrytime="00:00:32.84" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Salvador" lastname="Faustino" birthdate="1968-08-31" gender="M" nation="POR" license="119678" swrid="4610225" athleteid="42718">
              <RESULTS>
                <RESULT eventid="2537" points="322" reactiontime="+121" swimtime="00:01:36.05" resultid="42719" heatid="44886" lane="3" entrytime="00:01:33.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="331" reactiontime="+83" swimtime="00:00:39.93" resultid="42720" heatid="44896" lane="1" entrytime="00:00:36.84" />
                <RESULT eventid="2218" points="318" reactiontime="+86" swimtime="00:03:37.10" resultid="42721" heatid="44919" lane="8" entrytime="00:03:26.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.38" />
                    <SPLIT distance="100" swimtime="00:01:45.94" />
                    <SPLIT distance="150" swimtime="00:02:43.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="389" reactiontime="+81" swimtime="00:00:40.75" resultid="42722" heatid="45018" lane="3" entrytime="00:00:41.87" />
                <RESULT eventid="2652" points="419" reactiontime="+86" swimtime="00:00:33.57" resultid="42723" heatid="45041" lane="7" entrytime="00:00:31.24" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hugo Alexandre" lastname="Amaral" birthdate="1987-03-30" gender="M" nation="POR" license="12641" swrid="4064571" athleteid="42708">
              <RESULTS>
                <RESULT eventid="2682" points="555" reactiontime="+102" swimtime="00:00:30.43" resultid="42709" heatid="44897" lane="4" entrytime="00:00:32.67" />
                <RESULT eventid="2188" points="559" reactiontime="+79" swimtime="00:00:34.94" resultid="42710" heatid="44950" lane="8" entrytime="00:00:35.02" />
                <RESULT eventid="2445" points="449" reactiontime="+87" swimtime="00:01:23.39" resultid="42711" heatid="44998" lane="6" entrytime="00:01:20.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Andre" lastname="Mendonca" birthdate="1980-01-24" gender="M" nation="POR" license="25707" swrid="5003463" athleteid="42728">
              <RESULTS>
                <RESULT eventid="2652" points="607" reactiontime="+75" swimtime="00:00:29.03" resultid="42729" heatid="45045" lane="1" entrytime="00:00:28.44" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filipa Nobre" lastname="Chaveca" birthdate="1974-06-25" gender="F" nation="POR" license="210741" swrid="5376443" athleteid="42712">
              <RESULTS>
                <RESULT eventid="2203" points="241" reactiontime="+80" swimtime="00:01:53.02" resultid="42713" heatid="44881" lane="5" entrytime="00:01:46.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2278" points="225" reactiontime="+104" swimtime="00:03:39.03" resultid="42714" heatid="44903" lane="1" entrytime="00:03:20.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.36" />
                    <SPLIT distance="100" swimtime="00:01:44.33" />
                    <SPLIT distance="150" swimtime="00:02:43.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="280" reactiontime="+101" swimtime="00:01:31.58" resultid="42715" heatid="44953" lane="4" entrytime="00:01:36.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="221" reactiontime="+111" swimtime="00:00:51.81" resultid="42716" heatid="45024" lane="5" entrytime="00:00:50.99" entrycourse="LCM" />
                <RESULT eventid="2430" points="325" reactiontime="+113" swimtime="00:00:40.39" resultid="42717" heatid="45068" lane="7" entrytime="00:00:42.29" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara Andreia" lastname="Martins" birthdate="1981-11-03" gender="F" nation="POR" license="214295" athleteid="42724">
              <RESULTS>
                <RESULT eventid="2607" points="351" reactiontime="+102" swimtime="00:00:49.53" resultid="42725" heatid="45101" lane="7" entrytime="00:00:46.85" />
                <RESULT eventid="2522" points="217" reactiontime="+88" swimtime="00:00:52.70" resultid="42726" heatid="45025" lane="7" entrytime="00:00:45.97" />
                <RESULT eventid="2430" points="283" reactiontime="+100" swimtime="00:00:41.81" resultid="42727" heatid="45068" lane="5" entrytime="00:00:39.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ines Isabel" lastname="Silva" birthdate="1978-12-22" gender="F" nation="POR" license="103617" swrid="4660951" athleteid="42730">
              <RESULTS>
                <RESULT eventid="2338" points="397" reactiontime="+84" swimtime="00:00:39.93" resultid="42731" heatid="44891" lane="1" entrytime="00:00:37.93" entrycourse="SCM" />
                <RESULT eventid="2607" points="580" reactiontime="+83" swimtime="00:00:41.91" resultid="42732" heatid="45102" lane="7" entrytime="00:00:43.95" entrycourse="LCM" />
                <RESULT eventid="2460" points="507" reactiontime="+86" swimtime="00:01:36.32" resultid="42733" heatid="45121" lane="4" entrytime="00:01:40.87">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="531" reactiontime="+86" swimtime="00:00:33.88" resultid="42734" heatid="45071" lane="7" entrytime="00:00:33.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="VSC" nation="POR" region="ANNP" clubid="41926" swrid="65811" name="Vitoria Sport Clube" shortname="Vitoria Guimaraes">
          <ATHLETES>
            <ATHLETE firstname="David Nunes" lastname="Sousa" birthdate="1996-07-30" gender="M" nation="POR" license="112204" swrid="4411746" athleteid="43736">
              <RESULTS>
                <RESULT eventid="2507" status="WDR" swimtime="00:00:00.00" resultid="43737" entrytime="00:02:23.00" />
                <RESULT eventid="2385" status="WDR" swimtime="00:00:00.00" resultid="43738" entrytime="00:02:50.00" />
                <RESULT eventid="2445" status="WDR" swimtime="00:00:00.00" resultid="43739" entrytime="00:01:28.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edgar Manuel" lastname="Guimaraes" birthdate="1980-09-10" gender="M" nation="POR" license="110317" swrid="4372958" athleteid="43686">
              <RESULTS>
                <RESULT eventid="2188" points="413" reactiontime="+84" swimtime="00:00:40.94" resultid="43687" heatid="44940" lane="4" entrytime="00:00:50.00" entrycourse="LCM" />
                <RESULT eventid="2652" points="402" reactiontime="+82" swimtime="00:00:33.28" resultid="43688" heatid="45035" lane="6" entrytime="00:00:40.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agostinho Jorge" lastname="Sousa" birthdate="1981-09-21" gender="M" nation="POR" license="203962" swrid="5125755" athleteid="43732">
              <RESULTS>
                <RESULT eventid="2188" points="289" reactiontime="+97" swimtime="00:00:46.10" resultid="43733" heatid="44941" lane="8" entrytime="00:00:50.00" />
                <RESULT eventid="2652" points="339" reactiontime="+89" swimtime="00:00:35.22" resultid="43734" heatid="45034" lane="5" entrytime="00:00:43.00" />
                <RESULT eventid="2293" status="DNS" swimtime="00:00:00.00" resultid="43735" heatid="45017" lane="1" entrytime="00:00:48.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Renato Augusto" lastname="Oliveira" birthdate="1985-07-02" gender="M" nation="POR" license="124863" swrid="4005155" athleteid="43717">
              <RESULTS>
                <RESULT eventid="2682" points="212" reactiontime="+85" swimtime="00:00:42.74" resultid="43718" heatid="44894" lane="6" entrytime="00:00:43.08" entrycourse="LCM" />
                <RESULT eventid="2323" points="159" reactiontime="+93" swimtime="00:01:47.42" resultid="43719" heatid="44926" lane="7" entrytime="00:01:52.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="337" reactiontime="+87" swimtime="00:01:14.69" resultid="43720" heatid="45109" lane="2" entrytime="00:01:15.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="George Luiz" lastname="Junior" birthdate="1977-12-07" gender="M" nation="POR" license="214252" athleteid="43692">
              <RESULTS>
                <RESULT eventid="1058" points="274" swimtime="00:13:29.86" resultid="43693" heatid="45082" lane="8" entrytime="00:14:00.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.86" />
                    <SPLIT distance="200" swimtime="00:03:13.24" />
                    <SPLIT distance="300" swimtime="00:04:57.43" />
                    <SPLIT distance="400" swimtime="00:06:41.52" />
                    <SPLIT distance="500" swimtime="00:08:26.70" />
                    <SPLIT distance="600" swimtime="00:10:10.38" />
                    <SPLIT distance="700" swimtime="00:11:54.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="156" reactiontime="+118" swimtime="00:00:48.10" resultid="43694" heatid="44894" lane="2" entrytime="00:00:45.00" />
                <RESULT eventid="2507" points="245" reactiontime="+117" swimtime="00:03:09.21" resultid="43695" heatid="45092" lane="6" entrytime="00:03:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                    <SPLIT distance="100" swimtime="00:01:26.52" />
                    <SPLIT distance="150" swimtime="00:02:18.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="149" reactiontime="+115" swimtime="00:04:09.25" resultid="43696" heatid="44977" lane="6" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.50" />
                    <SPLIT distance="100" swimtime="00:01:56.43" />
                    <SPLIT distance="150" swimtime="00:03:19.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="264" reactiontime="+139" swimtime="00:06:36.15" resultid="43697" heatid="45126" lane="5" entrytime="00:07:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.70" />
                    <SPLIT distance="100" swimtime="00:01:28.70" />
                    <SPLIT distance="150" swimtime="00:02:19.02" />
                    <SPLIT distance="200" swimtime="00:03:10.24" />
                    <SPLIT distance="250" swimtime="00:04:02.39" />
                    <SPLIT distance="300" swimtime="00:04:54.98" />
                    <SPLIT distance="350" swimtime="00:05:47.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Manuel" lastname="Gomes" birthdate="1988-04-02" gender="M" nation="POR" license="16043" swrid="4559115" athleteid="43683">
              <RESULTS>
                <RESULT eventid="2622" points="519" reactiontime="+89" swimtime="00:02:58.54" resultid="43684" heatid="44879" lane="3" entrytime="00:02:45.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                    <SPLIT distance="100" swimtime="00:01:24.12" />
                    <SPLIT distance="150" swimtime="00:02:11.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="627" reactiontime="+80" swimtime="00:00:33.63" resultid="43685" heatid="44950" lane="3" entrytime="00:00:33.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nelson da Costa" lastname="Ramalhoto" birthdate="1969-06-13" gender="M" nation="POR" license="110369" swrid="4372974" athleteid="43727">
              <RESULTS>
                <RESULT eventid="2188" points="248" reactiontime="+103" swimtime="00:00:49.53" resultid="43728" heatid="44941" lane="3" entrytime="00:00:48.09" entrycourse="LCM" />
                <RESULT eventid="2415" points="223" reactiontime="+93" swimtime="00:01:33.67" resultid="43729" heatid="45105" lane="1" entrytime="00:01:34.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="277" reactiontime="+94" swimtime="00:01:51.13" resultid="43730" heatid="44993" lane="8" entrytime="00:01:52.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="244" reactiontime="+92" swimtime="00:00:40.17" resultid="43731" heatid="45035" lane="4" entrytime="00:00:39.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Armindo Manuel" lastname="Lobo" birthdate="1984-04-17" gender="M" nation="POR" license="118906" swrid="4590317" athleteid="43698">
              <RESULTS>
                <RESULT eventid="2682" points="472" reactiontime="+70" swimtime="00:00:32.77" resultid="43699" heatid="44897" lane="7" entrytime="00:00:34.80" entrycourse="LCM" />
                <RESULT eventid="2415" points="490" reactiontime="+70" swimtime="00:01:05.90" resultid="43700" heatid="45113" lane="6" entrytime="00:01:03.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="527" reactiontime="+78" swimtime="00:00:29.13" resultid="43701" heatid="45043" lane="6" entrytime="00:00:29.03" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Norberto Matos" lastname="Pereira" birthdate="1975-10-18" gender="M" nation="POR" license="111733" swrid="4403592" athleteid="43721">
              <RESULTS>
                <RESULT eventid="1058" points="243" swimtime="00:14:08.44" resultid="43722" heatid="45081" lane="2" entrytime="00:14:36.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.74" />
                    <SPLIT distance="200" swimtime="00:03:18.94" />
                    <SPLIT distance="300" swimtime="00:05:08.19" />
                    <SPLIT distance="400" swimtime="00:06:58.30" />
                    <SPLIT distance="500" swimtime="00:08:48.47" />
                    <SPLIT distance="600" swimtime="00:10:38.18" />
                    <SPLIT distance="700" swimtime="00:12:26.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2323" points="135" reactiontime="+93" swimtime="00:01:57.64" resultid="43723" heatid="44925" lane="4" entrytime="00:01:58.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="331" reactiontime="+99" swimtime="00:01:20.73" resultid="43724" heatid="45107" lane="2" entrytime="00:01:22.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="332" reactiontime="+91" swimtime="00:00:35.90" resultid="43725" heatid="45037" lane="7" entrytime="00:00:36.13" entrycourse="LCM" />
                <RESULT eventid="2248" points="194" reactiontime="+102" swimtime="00:08:42.39" resultid="43726" heatid="45058" lane="4" entrytime="00:08:50.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.83" />
                    <SPLIT distance="100" swimtime="00:02:02.00" />
                    <SPLIT distance="150" swimtime="00:03:21.87" />
                    <SPLIT distance="200" swimtime="00:04:38.44" />
                    <SPLIT distance="250" swimtime="00:05:47.62" />
                    <SPLIT distance="300" swimtime="00:06:59.74" />
                    <SPLIT distance="350" swimtime="00:07:52.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Catarina" lastname="Milhazes" birthdate="1985-11-17" gender="F" nation="POR" license="119706" swrid="4610246" athleteid="43707">
              <RESULTS>
                <RESULT eventid="2203" points="214" reactiontime="+83" swimtime="00:01:56.43" resultid="43708" heatid="44882" lane="8" entrytime="00:01:42.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2308" points="198" reactiontime="+87" swimtime="00:04:15.12" resultid="43709" heatid="44914" lane="5" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.86" />
                    <SPLIT distance="100" swimtime="00:02:03.55" />
                    <SPLIT distance="150" swimtime="00:03:09.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="196" reactiontime="+93" swimtime="00:00:56.17" resultid="43710" heatid="45099" lane="5" entrytime="00:00:51.36" entrycourse="LCM" />
                <RESULT eventid="2460" points="158" reactiontime="+83" swimtime="00:02:14.10" resultid="43711" heatid="45120" lane="4" entrytime="00:01:50.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Miguel" lastname="Bras" birthdate="1991-07-29" gender="M" nation="POR" license="23964" swrid="4559859" athleteid="43672">
              <RESULTS>
                <RESULT eventid="2507" points="447" reactiontime="+68" swimtime="00:02:31.30" resultid="43673" heatid="45095" lane="8" entrytime="00:02:27.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                    <SPLIT distance="100" swimtime="00:01:10.98" />
                    <SPLIT distance="150" swimtime="00:01:52.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="517" reactiontime="+70" swimtime="00:01:03.32" resultid="43674" heatid="45114" lane="2" entrytime="00:01:02.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="435" reactiontime="+68" swimtime="00:02:53.65" resultid="43675" heatid="44980" lane="3" entrytime="00:02:49.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                    <SPLIT distance="100" swimtime="00:01:23.89" />
                    <SPLIT distance="150" swimtime="00:02:15.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="552" reactiontime="+68" swimtime="00:00:28.34" resultid="43676" heatid="45046" lane="7" entrytime="00:00:27.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Miguel" lastname="Matos" birthdate="1992-06-09" gender="M" nation="POR" license="204167" swrid="4637824" athleteid="43702">
              <RESULTS>
                <RESULT eventid="2682" points="361" reactiontime="+103" swimtime="00:00:35.19" resultid="43703" heatid="44896" lane="2" entrytime="00:00:36.47" entrycourse="LCM" />
                <RESULT eventid="2415" points="373" reactiontime="+86" swimtime="00:01:11.79" resultid="43704" heatid="45110" lane="7" entrytime="00:01:12.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="401" reactiontime="+91" swimtime="00:05:40.17" resultid="43705" heatid="45128" lane="5" entrytime="00:06:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                    <SPLIT distance="100" swimtime="00:01:17.81" />
                    <SPLIT distance="150" swimtime="00:02:00.89" />
                    <SPLIT distance="200" swimtime="00:02:44.52" />
                    <SPLIT distance="250" swimtime="00:03:28.77" />
                    <SPLIT distance="300" swimtime="00:04:13.87" />
                    <SPLIT distance="350" swimtime="00:04:58.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="368" reactiontime="+80" swimtime="00:00:32.30" resultid="43706" heatid="45039" lane="4" entrytime="00:00:32.91" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Sofia" lastname="Alves" birthdate="1995-02-24" gender="F" nation="POR" license="25757" swrid="4561549" athleteid="43666">
              <RESULTS>
                <RESULT eventid="2278" points="740" reactiontime="+84" swimtime="00:02:21.21" resultid="43667" heatid="44905" lane="5" entrytime="00:02:19.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="100" swimtime="00:01:07.52" />
                    <SPLIT distance="150" swimtime="00:01:44.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="734" reactiontime="+76" swimtime="00:01:03.45" resultid="43668" heatid="44957" lane="6" entrytime="00:01:07.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="661" reactiontime="+77" swimtime="00:00:29.95" resultid="43669" heatid="45072" lane="3" entrytime="00:00:30.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marco Paulo" lastname="Azevedo" birthdate="1970-01-14" gender="M" nation="POR" license="214234" athleteid="43670">
              <RESULTS>
                <RESULT eventid="2652" points="345" reactiontime="+112" swimtime="00:00:35.79" resultid="43671" heatid="45034" lane="1" entrytime="00:00:45.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Orlando" lastname="Novais" birthdate="1978-10-20" gender="M" nation="POR" license="110370" swrid="4372968" athleteid="43712">
              <RESULTS>
                <RESULT eventid="2622" points="377" reactiontime="+91" swimtime="00:03:28.77" resultid="43713" heatid="44877" lane="6" entrytime="00:03:19.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.63" />
                    <SPLIT distance="100" swimtime="00:01:38.68" />
                    <SPLIT distance="150" swimtime="00:02:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="369" reactiontime="+92" swimtime="00:00:42.51" resultid="43714" heatid="44946" lane="6" entrytime="00:00:40.79" entrycourse="LCM" />
                <RESULT eventid="2445" points="346" reactiontime="+91" swimtime="00:01:37.74" resultid="43715" heatid="44996" lane="3" entrytime="00:01:31.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="286" reactiontime="+87" swimtime="00:00:37.29" resultid="43716" heatid="45038" lane="7" entrytime="00:00:34.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hamilton Kenji" lastname="Ida" birthdate="1973-11-11" gender="M" nation="BRA" license="212656" swrid="5425460" athleteid="43689">
              <RESULTS>
                <RESULT eventid="2507" points="364" reactiontime="+83" swimtime="00:02:47.09" resultid="43690" heatid="45092" lane="2" entrytime="00:03:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                    <SPLIT distance="100" swimtime="00:01:18.25" />
                    <SPLIT distance="150" swimtime="00:02:02.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="382" reactiontime="+89" swimtime="00:05:52.96" resultid="43691" heatid="45126" lane="3" entrytime="00:07:00.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                    <SPLIT distance="100" swimtime="00:01:20.53" />
                    <SPLIT distance="150" swimtime="00:02:04.19" />
                    <SPLIT distance="200" swimtime="00:02:49.82" />
                    <SPLIT distance="250" swimtime="00:03:35.87" />
                    <SPLIT distance="300" swimtime="00:04:22.85" />
                    <SPLIT distance="350" swimtime="00:05:08.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Manuela" lastname="Ferreira" birthdate="1970-07-16" gender="F" nation="POR" license="130114" swrid="4988912" athleteid="43677">
              <RESULTS>
                <RESULT eventid="1060" points="271" swimtime="00:15:15.02" resultid="43678" heatid="45076" lane="4" entrytime="00:14:24.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.72" />
                    <SPLIT distance="200" swimtime="00:03:30.92" />
                    <SPLIT distance="300" swimtime="00:05:27.88" />
                    <SPLIT distance="400" swimtime="00:07:27.27" />
                    <SPLIT distance="500" swimtime="00:09:27.24" />
                    <SPLIT distance="600" swimtime="00:11:24.73" />
                    <SPLIT distance="700" swimtime="00:13:30.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2278" points="305" reactiontime="+90" swimtime="00:03:25.14" resultid="43679" heatid="44903" lane="7" entrytime="00:03:20.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.21" />
                    <SPLIT distance="100" swimtime="00:01:35.57" />
                    <SPLIT distance="150" swimtime="00:02:30.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="235" reactiontime="+113" swimtime="00:04:15.69" resultid="43680" heatid="44971" lane="4" entrytime="00:04:06.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.78" />
                    <SPLIT distance="100" swimtime="00:02:12.42" />
                    <SPLIT distance="150" swimtime="00:03:24.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="276" reactiontime="+104" swimtime="00:07:22.74" resultid="43681" heatid="45011" lane="1" entrytime="00:06:56.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.91" />
                    <SPLIT distance="100" swimtime="00:01:42.91" />
                    <SPLIT distance="150" swimtime="00:02:38.82" />
                    <SPLIT distance="200" swimtime="00:03:36.07" />
                    <SPLIT distance="250" swimtime="00:04:32.51" />
                    <SPLIT distance="300" swimtime="00:05:30.06" />
                    <SPLIT distance="350" swimtime="00:06:27.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="352" reactiontime="+92" swimtime="00:00:40.22" resultid="43682" heatid="45067" lane="6" entrytime="00:00:45.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="FOCA" nation="POR" region="ANNP" clubid="42401" swrid="66457" name="Foca-Clube Natacao de Felgueiras" shortname="Foca Quinta da Lixa CNF">
          <ATHLETES>
            <ATHLETE firstname="Luis Manuel" lastname="Ribeiro" birthdate="1991-07-27" gender="M" nation="POR" license="107830" swrid="5326937" athleteid="42430">
              <RESULTS>
                <RESULT eventid="2507" points="487" reactiontime="+82" swimtime="00:02:27.00" resultid="42431" heatid="45093" lane="6" entrytime="00:02:46.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="100" swimtime="00:01:10.40" />
                    <SPLIT distance="150" swimtime="00:01:49.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="427" reactiontime="+77" swimtime="00:00:38.22" resultid="42432" heatid="44946" lane="1" entrytime="00:00:41.15" />
                <RESULT eventid="2415" points="525" reactiontime="+81" swimtime="00:01:02.99" resultid="42433" heatid="45112" lane="3" entrytime="00:01:05.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="411" reactiontime="+80" swimtime="00:01:25.93" resultid="42434" heatid="44996" lane="5" entrytime="00:01:30.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="571" reactiontime="+76" swimtime="00:00:28.01" resultid="42435" heatid="45044" lane="1" entrytime="00:00:28.88" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose" lastname="Leite" birthdate="1948-09-16" gender="M" nation="POR" license="204547" swrid="5207388" athleteid="42412">
              <RESULTS>
                <RESULT eventid="2622" points="411" reactiontime="+120" swimtime="00:04:18.95" resultid="42413" heatid="44874" lane="2" entrytime="00:04:11.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.44" />
                    <SPLIT distance="100" swimtime="00:02:06.23" />
                    <SPLIT distance="150" swimtime="00:03:15.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="356" reactiontime="+109" swimtime="00:00:51.99" resultid="42414" heatid="44940" lane="6" entrytime="00:00:50.61" />
                <RESULT eventid="2445" points="348" reactiontime="+109" swimtime="00:02:01.81" resultid="42415" heatid="44992" lane="5" entrytime="00:01:54.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Brandao" lastname="Andrade" birthdate="1949-06-24" gender="M" nation="POR" license="153287" swrid="5115761" athleteid="42402">
              <RESULTS>
                <RESULT eventid="2188" points="198" reactiontime="+135" swimtime="00:01:03.20" resultid="42403" heatid="44938" lane="4" entrytime="00:01:00.67" />
                <RESULT eventid="2652" points="65" reactiontime="+132" swimtime="00:01:10.77" resultid="42404" heatid="45032" lane="4" entrytime="00:01:01.33" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mario Nuno" lastname="Pereira" birthdate="1981-02-20" gender="M" nation="POR" license="200652" swrid="5157491" athleteid="42423">
              <RESULTS>
                <RESULT eventid="2263" points="306" reactiontime="+107" swimtime="00:06:17.09" resultid="42424" heatid="45128" lane="1" entrytime="00:06:28.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                    <SPLIT distance="100" swimtime="00:01:25.55" />
                    <SPLIT distance="150" swimtime="00:02:12.60" />
                    <SPLIT distance="200" swimtime="00:03:02.04" />
                    <SPLIT distance="250" swimtime="00:03:50.45" />
                    <SPLIT distance="300" swimtime="00:04:40.55" />
                    <SPLIT distance="350" swimtime="00:05:30.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="42425" heatid="45039" lane="3" entrytime="00:00:33.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filipe Pinheiro" lastname="Pires" birthdate="1973-05-02" gender="M" nation="POR" license="117638" swrid="4557827" athleteid="42426">
              <RESULTS>
                <RESULT eventid="1058" points="355" swimtime="00:12:28.53" resultid="42427" heatid="45083" lane="6" entrytime="00:12:39.03">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.73" />
                    <SPLIT distance="200" swimtime="00:03:00.07" />
                    <SPLIT distance="300" swimtime="00:04:34.32" />
                    <SPLIT distance="400" swimtime="00:06:10.29" />
                    <SPLIT distance="500" swimtime="00:07:45.64" />
                    <SPLIT distance="600" swimtime="00:09:21.36" />
                    <SPLIT distance="700" swimtime="00:10:56.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" status="DNS" swimtime="00:00:00.00" resultid="42428" heatid="45128" lane="2" entrytime="00:06:15.61" />
                <RESULT eventid="2415" points="393" reactiontime="+88" swimtime="00:01:16.23" resultid="42429" heatid="45105" lane="2" entrytime="00:01:32.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor Carvalho" lastname="Lopes" birthdate="1972-09-24" gender="M" nation="POR" license="132421" swrid="5068135" athleteid="42416">
              <RESULTS>
                <RESULT eventid="2188" points="305" reactiontime="+106" swimtime="00:00:44.41" resultid="42417" heatid="44945" lane="2" entrytime="00:00:42.69" />
                <RESULT eventid="2445" points="330" reactiontime="+101" swimtime="00:01:39.64" resultid="42418" heatid="44996" lane="1" entrytime="00:01:34.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Albano Couto" lastname="Teixeira" birthdate="1963-08-30" gender="M" nation="POR" license="117114" swrid="5068174" athleteid="42436">
              <RESULTS>
                <RESULT eventid="2622" points="247" reactiontime="+115" swimtime="00:04:20.21" resultid="42437" heatid="44873" lane="3" entrytime="00:04:27.94">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.71" />
                    <SPLIT distance="100" swimtime="00:02:00.77" />
                    <SPLIT distance="150" swimtime="00:03:10.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="197" reactiontime="+117" swimtime="00:00:53.33" resultid="42438" heatid="44940" lane="1" entrytime="00:00:51.36" />
                <RESULT comment="733 - Efectuou varias braçadas durante percurso subaquático após a partida - SW 7.1" eventid="2445" reactiontime="+115" status="DSQ" swimtime="00:01:58.49" resultid="42439" heatid="44992" lane="1" entrytime="00:01:59.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rosa Leitao" lastname="Costa" birthdate="1965-07-15" gender="F" nation="POR" license="132419" swrid="5068113" athleteid="42405">
              <RESULTS>
                <RESULT eventid="2607" points="282" reactiontime="+110" swimtime="00:00:57.61" resultid="42406" heatid="45098" lane="6" entrytime="00:00:58.52" />
                <RESULT eventid="2460" points="323" reactiontime="+110" swimtime="00:02:03.48" resultid="42407" heatid="45119" lane="2" entrytime="00:02:02.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2173" points="403" swimtime="00:04:16.28" resultid="42408" heatid="45087" lane="6" entrytime="00:04:15.54">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.79" />
                    <SPLIT distance="100" swimtime="00:02:01.67" />
                    <SPLIT distance="150" swimtime="00:03:09.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuel Fernando" lastname="Fernandes" birthdate="1968-03-14" gender="M" nation="POR" license="202748" swrid="4845987" athleteid="42409">
              <RESULTS>
                <RESULT eventid="2445" points="222" reactiontime="+117" swimtime="00:01:59.58" resultid="42410" heatid="44991" lane="4" entrytime="00:02:02.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="208" reactiontime="+111" swimtime="00:00:52.54" resultid="42411" heatid="44939" lane="5" entrytime="00:00:52.16" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raquel Filipa" lastname="Miranda" birthdate="1985-02-03" gender="F" nation="POR" license="132422" swrid="4564416" athleteid="42419">
              <RESULTS>
                <RESULT eventid="2203" points="542" reactiontime="+102" swimtime="00:01:25.45" resultid="42420" heatid="44883" lane="2" entrytime="00:01:23.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="608" reactiontime="+95" swimtime="00:02:56.07" resultid="42421" heatid="44974" lane="2" entrytime="00:02:55.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.72" />
                    <SPLIT distance="100" swimtime="00:01:27.02" />
                    <SPLIT distance="150" swimtime="00:02:16.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="441" reactiontime="+87" swimtime="00:01:35.31" resultid="42422" heatid="45123" lane="7" entrytime="00:01:30.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CDE" nation="POR" region="ANCNP" clubid="41800" swrid="68060" name="Clube Desportivo Estarreja" shortname="Estarreja">
          <ATHLETES>
            <ATHLETE firstname="Olivia Cristina" lastname="Nunes" birthdate="1972-06-02" gender="F" nation="POR" license="209367" swrid="5336583" athleteid="41812">
              <RESULTS>
                <RESULT eventid="2173" points="145" swimtime="00:05:24.68" resultid="41813" heatid="45086" lane="5" entrytime="00:05:01.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.00" />
                    <SPLIT distance="100" swimtime="00:02:35.68" />
                    <SPLIT distance="150" swimtime="00:04:02.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2338" points="96" reactiontime="+151" swimtime="00:01:05.88" resultid="41814" heatid="44889" lane="2" entrytime="00:01:05.00" />
                <RESULT eventid="2607" points="162" reactiontime="+130" swimtime="00:01:06.38" resultid="41815" heatid="45098" lane="1" entrytime="00:01:02.67" entrycourse="LCM" />
                <RESULT eventid="2460" points="161" reactiontime="+130" swimtime="00:02:27.13" resultid="41816" heatid="45118" lane="5" entrytime="00:02:20.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="111" reactiontime="+122" swimtime="00:00:57.75" resultid="41817" heatid="45066" lane="6" entrytime="00:00:54.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Renato Castro" lastname="Valente" birthdate="1979-10-30" gender="M" nation="POR" license="209675" swrid="5344117" athleteid="41835">
              <RESULTS>
                <RESULT eventid="2537" points="332" reactiontime="+99" swimtime="00:01:28.58" resultid="41836" heatid="44887" lane="8" entrytime="00:01:31.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="376" reactiontime="+92" swimtime="00:00:42.25" resultid="41837" heatid="44946" lane="8" entrytime="00:00:41.84" entrycourse="LCM" />
                <RESULT eventid="2415" points="396" reactiontime="+95" swimtime="00:01:13.97" resultid="41838" heatid="45110" lane="8" entrytime="00:01:13.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="400" reactiontime="+67" swimtime="00:00:38.54" resultid="41839" heatid="45018" lane="4" entrytime="00:00:40.95" entrycourse="LCM" />
                <RESULT eventid="2652" points="512" reactiontime="+92" swimtime="00:00:30.72" resultid="41840" heatid="45040" lane="3" entrytime="00:00:31.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago Sousa" lastname="Tavares" birthdate="1984-09-23" gender="M" nation="POR" license="108108" swrid="4319442" athleteid="41827">
              <RESULTS>
                <RESULT eventid="1058" status="DNS" swimtime="00:00:00.00" resultid="41828" heatid="45083" lane="3" entrytime="00:12:30.00" />
                <RESULT eventid="2507" status="DNS" swimtime="00:00:00.00" resultid="41829" heatid="45094" lane="5" entrytime="00:02:29.80" />
                <RESULT eventid="2385" status="DNS" swimtime="00:00:00.00" resultid="41830" heatid="44980" lane="8" entrytime="00:02:55.00" />
                <RESULT eventid="2263" status="DNS" swimtime="00:00:00.00" resultid="41831" heatid="45129" lane="4" entrytime="00:05:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel Angelo" lastname="Nunes" birthdate="1973-05-31" gender="M" nation="POR" license="206646" swrid="5278981" athleteid="41806">
              <RESULTS>
                <RESULT eventid="2622" points="467" reactiontime="+83" swimtime="00:03:18.06" resultid="41807" heatid="44877" lane="1" entrytime="00:03:20.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.76" />
                    <SPLIT distance="100" swimtime="00:01:33.22" />
                    <SPLIT distance="150" swimtime="00:02:25.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="463" reactiontime="+81" swimtime="00:00:34.32" resultid="41808" heatid="44897" lane="6" entrytime="00:00:34.03" entrycourse="LCM" />
                <RESULT eventid="2188" points="420" reactiontime="+78" swimtime="00:00:39.90" resultid="41809" heatid="44947" lane="2" entrytime="00:00:39.07" entrycourse="LCM" />
                <RESULT eventid="2385" points="465" reactiontime="+85" swimtime="00:02:57.67" resultid="41810" heatid="44979" lane="4" entrytime="00:02:55.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:24.09" />
                    <SPLIT distance="150" swimtime="00:02:17.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="441" reactiontime="+84" swimtime="00:06:37.25" resultid="41811" heatid="45061" lane="6" entrytime="00:06:21.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                    <SPLIT distance="100" swimtime="00:01:25.53" />
                    <SPLIT distance="150" swimtime="00:02:20.83" />
                    <SPLIT distance="200" swimtime="00:03:15.74" />
                    <SPLIT distance="250" swimtime="00:04:13.73" />
                    <SPLIT distance="300" swimtime="00:05:11.41" />
                    <SPLIT distance="350" swimtime="00:05:55.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Pedro" lastname="Santos" birthdate="1995-06-17" gender="M" nation="POR" license="105859" swrid="4251289" athleteid="41823">
              <RESULTS>
                <RESULT eventid="2415" points="769" reactiontime="+68" swimtime="00:00:56.43" resultid="41824" heatid="45116" lane="1" entrytime="00:00:57.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="792" reactiontime="+83" swimtime="00:00:28.94" resultid="41825" heatid="45022" lane="5" entrytime="00:00:30.00" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="41826" heatid="45047" lane="1" entrytime="00:00:27.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Elisabete" lastname="Oliveira" birthdate="1949-03-25" gender="F" nation="POR" license="211854" swrid="5425458" athleteid="41818">
              <RESULTS>
                <RESULT eventid="2607" points="114" swimtime="00:01:25.81" resultid="41819" heatid="45097" lane="1" entrytime="00:02:00.00" />
                <RESULT eventid="2460" points="127" swimtime="00:03:21.07" resultid="41820" heatid="45118" lane="1" entrytime="00:03:50.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:33.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2522" points="115" reactiontime="+86" swimtime="00:01:26.98" resultid="41821" heatid="45023" lane="8" entrytime="00:01:45.00" />
                <RESULT eventid="2430" points="109" swimtime="00:01:10.08" resultid="41822" heatid="45065" lane="5" entrytime="00:01:10.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nuno Ricardo" lastname="Ferreira" birthdate="1985-10-22" gender="M" nation="POR" license="213021" swrid="5447637" athleteid="41801">
              <RESULTS>
                <RESULT eventid="2188" points="148" reactiontime="+101" swimtime="00:00:55.10" resultid="41802" heatid="44940" lane="8" entrytime="00:00:51.68" entrycourse="LCM" />
                <RESULT eventid="2415" points="139" reactiontime="+96" swimtime="00:01:40.27" resultid="41803" heatid="45104" lane="3" entrytime="00:01:45.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="156" reactiontime="+94" swimtime="00:02:03.33" resultid="41804" heatid="44992" lane="8" entrytime="00:02:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="172" reactiontime="+84" swimtime="00:00:42.31" resultid="41805" heatid="45034" lane="3" entrytime="00:00:43.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre Manuel" lastname="Teixeira" birthdate="1978-07-21" gender="M" nation="POR" license="208841" swrid="5330800" athleteid="41832">
              <RESULTS>
                <RESULT eventid="2188" points="247" reactiontime="+86" swimtime="00:00:48.62" resultid="41833" heatid="44942" lane="8" entrytime="00:00:47.14" entrycourse="LCM" />
                <RESULT eventid="2385" points="255" reactiontime="+89" swimtime="00:03:28.64" resultid="41834" heatid="44977" lane="4" entrytime="00:03:15.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:01:33.75" />
                    <SPLIT distance="150" swimtime="00:02:37.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="ACS" nation="POR" region="ANALG" clubid="43061" swrid="84075" name="Aquatico Clube de Silves" shortname="Aquatico Silves">
          <ATHLETES>
            <ATHLETE firstname="Joana Isabel" lastname="Cunha" birthdate="1980-07-17" gender="F" nation="POR" license="117125" swrid="4475974" athleteid="43062">
              <RESULTS>
                <RESULT eventid="2607" points="584" reactiontime="+75" swimtime="00:00:41.82" resultid="43063" heatid="45103" lane="2" entrytime="00:00:40.50" />
                <RESULT eventid="2637" points="626" reactiontime="+70" swimtime="00:01:10.49" resultid="43064" heatid="44957" lane="8" entrytime="00:01:10.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="618" reactiontime="+69" swimtime="00:02:57.77" resultid="43065" heatid="44974" lane="7" entrytime="00:02:55.67">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:25.38" />
                    <SPLIT distance="150" swimtime="00:02:17.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="541" reactiontime="+73" swimtime="00:05:46.87" resultid="43066" heatid="45013" lane="6" entrytime="00:05:30.84">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                    <SPLIT distance="100" swimtime="00:01:17.22" />
                    <SPLIT distance="150" swimtime="00:02:01.37" />
                    <SPLIT distance="200" swimtime="00:02:45.93" />
                    <SPLIT distance="250" swimtime="00:03:31.55" />
                    <SPLIT distance="300" swimtime="00:04:17.33" />
                    <SPLIT distance="350" swimtime="00:05:03.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2400" points="618" reactiontime="+77" swimtime="00:06:20.78" resultid="43067" heatid="45064" lane="5" entrytime="00:06:05.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                    <SPLIT distance="100" swimtime="00:01:23.23" />
                    <SPLIT distance="150" swimtime="00:02:17.49" />
                    <SPLIT distance="200" swimtime="00:03:08.25" />
                    <SPLIT distance="250" swimtime="00:04:01.31" />
                    <SPLIT distance="300" swimtime="00:04:54.40" />
                    <SPLIT distance="350" swimtime="00:05:37.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CGA" nation="POR" region="ANCNP" clubid="41928" swrid="72840" name="Clube dos Galitos" shortname="Galitos/ Bresimar">
          <ATHLETES>
            <ATHLETE firstname="Nuno Alexandre" lastname="Lobo" birthdate="1970-10-01" gender="M" nation="POR" license="210712" swrid="5376438" athleteid="42487">
              <RESULTS>
                <RESULT eventid="2218" points="543" reactiontime="+72" swimtime="00:03:01.79" resultid="42488" heatid="44920" lane="2" entrytime="00:02:58.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                    <SPLIT distance="100" swimtime="00:01:25.27" />
                    <SPLIT distance="150" swimtime="00:02:16.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="578" reactiontime="+96" swimtime="00:00:37.36" resultid="42489" heatid="44949" lane="1" entrytime="00:00:36.10" />
                <RESULT eventid="2293" points="613" reactiontime="+70" swimtime="00:00:35.02" resultid="42490" heatid="45021" lane="7" entrytime="00:00:33.18" entrycourse="SCM" />
                <RESULT eventid="2652" points="726" reactiontime="+90" swimtime="00:00:27.94" resultid="42491" heatid="45045" lane="5" entrytime="00:00:27.86" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Rosas" lastname="Lobo" birthdate="1983-02-23" gender="M" nation="POR" license="148709" swrid="5106685" athleteid="42482">
              <RESULTS>
                <RESULT eventid="2682" points="706" reactiontime="+74" swimtime="00:00:28.65" resultid="42483" heatid="44901" lane="8" entrytime="00:00:28.53" entrycourse="LCM" />
                <RESULT eventid="2323" points="653" reactiontime="+84" swimtime="00:01:07.11" resultid="42484" heatid="44930" lane="7" entrytime="00:01:04.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="616" reactiontime="+79" swimtime="00:01:01.07" resultid="42485" heatid="45115" lane="3" entrytime="00:00:59.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="592" reactiontime="+80" swimtime="00:00:28.02" resultid="42486" heatid="45047" lane="5" entrytime="00:00:26.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo Ferreira" lastname="Basto" birthdate="1967-06-28" gender="M" nation="POR" license="103219" swrid="4607041" athleteid="42473">
              <RESULTS>
                <RESULT eventid="2622" points="551" reactiontime="+86" swimtime="00:03:15.13" resultid="42474" heatid="44878" lane="8" entrytime="00:03:17.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                    <SPLIT distance="100" swimtime="00:01:32.17" />
                    <SPLIT distance="150" swimtime="00:02:24.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2323" points="462" reactiontime="+85" swimtime="00:01:22.35" resultid="42475" heatid="44927" lane="6" entrytime="00:01:21.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="534" reactiontime="+87" swimtime="00:02:57.67" resultid="42476" heatid="44979" lane="3" entrytime="00:02:57.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="100" swimtime="00:01:22.72" />
                    <SPLIT distance="150" swimtime="00:02:14.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" points="406" reactiontime="+99" swimtime="00:03:18.62" resultid="42477" heatid="45029" lane="4" entrytime="00:03:15.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.12" />
                    <SPLIT distance="100" swimtime="00:01:35.69" />
                    <SPLIT distance="150" swimtime="00:02:30.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="521" reactiontime="+98" swimtime="00:06:34.24" resultid="42478" heatid="45060" lane="3" entrytime="00:06:35.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:01:26.26" />
                    <SPLIT distance="150" swimtime="00:02:18.61" />
                    <SPLIT distance="200" swimtime="00:03:11.17" />
                    <SPLIT distance="250" swimtime="00:04:06.43" />
                    <SPLIT distance="300" swimtime="00:05:03.10" />
                    <SPLIT distance="350" swimtime="00:05:50.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Celso Filipe" lastname="Assuncao" birthdate="1978-11-16" gender="M" nation="POR" license="125458" swrid="4405287" athleteid="42469">
              <RESULTS>
                <RESULT eventid="2188" points="677" reactiontime="+80" swimtime="00:00:34.74" resultid="42470" heatid="44950" lane="1" entrytime="00:00:34.34" entrycourse="LCM" />
                <RESULT eventid="2445" points="638" reactiontime="+75" swimtime="00:01:19.73" resultid="42471" heatid="44998" lane="2" entrytime="00:01:22.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="597" reactiontime="+73" swimtime="00:00:29.19" resultid="42472" heatid="45043" lane="2" entrytime="00:00:29.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Margarida" lastname="Rodrigues" birthdate="1996-09-03" gender="F" nation="POR" license="103868" swrid="4251302" athleteid="42498">
              <RESULTS>
                <RESULT eventid="2338" points="785" reactiontime="+78" swimtime="00:00:30.13" resultid="42499" heatid="44892" lane="4" entrytime="00:00:28.53" entrycourse="LCM" />
                <RESULT eventid="2278" points="734" reactiontime="+87" swimtime="00:02:21.62" resultid="42500" heatid="44905" lane="4" entrytime="00:02:10.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:07.83" />
                    <SPLIT distance="150" swimtime="00:01:45.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2552" points="739" reactiontime="+85" swimtime="00:01:08.67" resultid="42501" heatid="44924" lane="4" entrytime="00:01:02.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="730" reactiontime="+82" swimtime="00:02:38.30" resultid="42502" heatid="44974" lane="4" entrytime="00:02:29.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                    <SPLIT distance="100" swimtime="00:01:14.41" />
                    <SPLIT distance="150" swimtime="00:02:02.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" status="WDR" swimtime="00:00:00.00" resultid="42503" entrytime="00:00:28.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo Lourenco" lastname="Alves" birthdate="1984-05-02" gender="M" nation="POR" license="203281" swrid="4940915" athleteid="42466">
              <RESULTS>
                <RESULT eventid="1058" points="332" swimtime="00:12:53.36" resultid="42467" heatid="45083" lane="4" entrytime="00:12:14.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.01" />
                    <SPLIT distance="200" swimtime="00:02:59.33" />
                    <SPLIT distance="300" swimtime="00:04:37.36" />
                    <SPLIT distance="400" swimtime="00:06:17.09" />
                    <SPLIT distance="500" swimtime="00:07:58.69" />
                    <SPLIT distance="600" swimtime="00:09:38.14" />
                    <SPLIT distance="700" swimtime="00:11:17.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" status="WDR" swimtime="00:00:00.00" resultid="42468" entrytime="00:02:54.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Henrique" lastname="Madail" birthdate="1954-11-15" gender="M" nation="POR" license="119658" swrid="4607101" athleteid="42492">
              <RESULTS>
                <RESULT eventid="1058" points="287" swimtime="00:16:20.39" resultid="42493" heatid="45080" lane="5" entrytime="00:15:44.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.88" />
                    <SPLIT distance="200" swimtime="00:03:59.29" />
                    <SPLIT distance="300" swimtime="00:06:03.83" />
                    <SPLIT distance="400" swimtime="00:08:08.36" />
                    <SPLIT distance="500" swimtime="00:10:12.75" />
                    <SPLIT distance="600" swimtime="00:12:17.35" />
                    <SPLIT distance="700" swimtime="00:14:21.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="284" reactiontime="+89" swimtime="00:00:52.49" resultid="42494" heatid="44941" lane="1" entrytime="00:00:49.83" entrycourse="LCM" />
                <RESULT eventid="2263" points="315" reactiontime="+96" swimtime="00:07:41.81" resultid="42495" heatid="45125" lane="4" entrytime="00:07:43.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.97" />
                    <SPLIT distance="100" swimtime="00:01:44.85" />
                    <SPLIT distance="150" swimtime="00:02:44.22" />
                    <SPLIT distance="200" swimtime="00:03:45.48" />
                    <SPLIT distance="250" swimtime="00:04:46.02" />
                    <SPLIT distance="300" swimtime="00:05:46.86" />
                    <SPLIT distance="350" swimtime="00:06:46.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="381" reactiontime="+99" swimtime="00:01:53.62" resultid="42496" heatid="44992" lane="3" entrytime="00:01:55.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="42497" heatid="45034" lane="7" entrytime="00:00:44.89" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo Jorge" lastname="Jesus" birthdate="1975-06-21" gender="M" nation="POR" license="206044" swrid="5261138" athleteid="42479">
              <RESULTS>
                <RESULT eventid="2293" points="520" reactiontime="+104" swimtime="00:00:35.76" resultid="42480" heatid="45021" lane="1" entrytime="00:00:33.37" entrycourse="SCM" />
                <RESULT eventid="2652" points="609" reactiontime="+77" swimtime="00:00:29.33" resultid="42481" heatid="45044" lane="8" entrytime="00:00:28.92" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GAN" nation="POR" region="ANL" clubid="41726" swrid="85652" name="Grupo dos Amigos da Natacao-ACD" shortname="Amigos da Natacao">
          <ATHLETES>
            <ATHLETE firstname="Anabela Verissimo" lastname="Mota" birthdate="1966-04-23" gender="F" nation="POR" license="206914" swrid="5276376" athleteid="41754">
              <RESULTS>
                <RESULT eventid="1060" points="181" swimtime="00:17:47.80" resultid="41755" heatid="45074" lane="6" entrytime="00:18:15.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:05.85" />
                    <SPLIT distance="200" swimtime="00:04:20.18" />
                    <SPLIT distance="300" swimtime="00:06:33.46" />
                    <SPLIT distance="400" swimtime="00:08:48.05" />
                    <SPLIT distance="500" swimtime="00:11:01.70" />
                    <SPLIT distance="600" swimtime="00:13:18.06" />
                    <SPLIT distance="700" swimtime="00:15:36.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2338" points="148" reactiontime="+114" swimtime="00:01:00.17" resultid="41756" heatid="44889" lane="5" entrytime="00:00:59.33" entrycourse="LCM" />
                <RESULT comment="atleta a partir dos 20 metros mudou de estilo" eventid="2552" reactiontime="+113" status="DSQ" swimtime="00:02:28.76" resultid="41757" heatid="44922" lane="5" entrytime="00:02:09.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="197" reactiontime="+114" swimtime="00:01:49.42" resultid="41758" heatid="44953" lane="8" entrytime="00:01:51.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="283" reactiontime="+107" swimtime="00:00:45.10" resultid="41759" heatid="45067" lane="1" entrytime="00:00:46.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nuno Silva" lastname="Afonso" birthdate="1979-12-15" gender="M" nation="POR" license="201498" swrid="5171531" athleteid="41748">
              <RESULTS>
                <RESULT eventid="1058" points="217" swimtime="00:14:35.30" resultid="41749" heatid="45081" lane="4" entrytime="00:15:38.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.30" />
                    <SPLIT distance="200" swimtime="00:03:23.87" />
                    <SPLIT distance="300" swimtime="00:05:16.73" />
                    <SPLIT distance="400" swimtime="00:07:11.21" />
                    <SPLIT distance="500" swimtime="00:09:05.38" />
                    <SPLIT distance="600" swimtime="00:10:59.49" />
                    <SPLIT distance="700" swimtime="00:12:51.63" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="604 - Durante o percurso perdeu a posição dorsal - SW 6.2" eventid="2218" reactiontime="+76" status="DSQ" swimtime="00:03:48.66" resultid="41750" heatid="44920" lane="6" entrytime="00:03:57.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.33" />
                    <SPLIT distance="100" swimtime="00:01:51.56" />
                    <SPLIT distance="150" swimtime="00:02:50.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="243" reactiontime="+116" swimtime="00:03:32.15" resultid="41751" heatid="44977" lane="1" entrytime="00:03:35.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.62" />
                    <SPLIT distance="100" swimtime="00:01:47.58" />
                    <SPLIT distance="150" swimtime="00:02:44.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" points="163" reactiontime="+129" swimtime="00:04:02.07" resultid="41752" heatid="45029" lane="1" entrytime="00:04:00.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.30" />
                    <SPLIT distance="100" swimtime="00:01:55.61" />
                    <SPLIT distance="150" swimtime="00:03:00.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="303" reactiontime="+102" swimtime="00:00:36.57" resultid="41753" heatid="45034" lane="4" entrytime="00:00:42.86" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago Filipe" lastname="Cunha" birthdate="1976-05-07" gender="M" nation="POR" license="204756" swrid="5215228" athleteid="41736">
              <RESULTS>
                <RESULT eventid="2622" points="438" reactiontime="+89" swimtime="00:03:22.32" resultid="41737" heatid="44876" lane="2" entrytime="00:03:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.11" />
                    <SPLIT distance="100" swimtime="00:01:36.40" />
                    <SPLIT distance="150" swimtime="00:02:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="340" reactiontime="+88" swimtime="00:01:19.97" resultid="41738" heatid="45107" lane="7" entrytime="00:01:22.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="381" reactiontime="+97" swimtime="00:03:09.88" resultid="41739" heatid="44977" lane="5" entrytime="00:03:18.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.08" />
                    <SPLIT distance="100" swimtime="00:01:34.77" />
                    <SPLIT distance="150" swimtime="00:02:25.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="423" reactiontime="+88" swimtime="00:01:31.77" resultid="41740" heatid="44996" lane="7" entrytime="00:01:33.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="394" reactiontime="+91" swimtime="00:06:52.47" resultid="41741" heatid="45060" lane="8" entrytime="00:07:02.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                    <SPLIT distance="100" swimtime="00:01:38.17" />
                    <SPLIT distance="150" swimtime="00:02:33.13" />
                    <SPLIT distance="200" swimtime="00:03:26.17" />
                    <SPLIT distance="250" swimtime="00:04:21.93" />
                    <SPLIT distance="300" swimtime="00:05:18.16" />
                    <SPLIT distance="350" swimtime="00:06:06.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Pedro" lastname="Marques" birthdate="1977-10-23" gender="M" nation="POR" license="206630" swrid="5276374" athleteid="41727">
              <RESULTS>
                <RESULT eventid="2293" status="DNS" swimtime="00:00:00.00" resultid="41728" heatid="45014" lane="8" entrytime="00:01:15.00" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="41729" heatid="45038" lane="6" entrytime="00:00:34.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Maria" lastname="Caeiro" birthdate="1959-02-15" gender="F" nation="POR" license="201953" swrid="5191870" athleteid="41742">
              <RESULTS>
                <RESULT eventid="1060" points="364" swimtime="00:16:30.06" resultid="41743" heatid="45076" lane="1" entrytime="00:15:47.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.99" />
                    <SPLIT distance="200" swimtime="00:04:01.07" />
                    <SPLIT distance="300" swimtime="00:06:07.45" />
                    <SPLIT distance="400" swimtime="00:08:13.19" />
                    <SPLIT distance="500" swimtime="00:10:19.01" />
                    <SPLIT distance="600" swimtime="00:12:24.58" />
                    <SPLIT distance="700" swimtime="00:14:29.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2338" points="176" reactiontime="+121" swimtime="00:00:59.55" resultid="41744" heatid="44890" lane="8" entrytime="00:00:54.54" entrycourse="LCM" />
                <RESULT eventid="2552" points="220" reactiontime="+129" swimtime="00:02:14.44" resultid="41745" heatid="44922" lane="3" entrytime="00:02:09.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="261" reactiontime="+129" swimtime="00:04:38.40" resultid="41746" heatid="44971" lane="2" entrytime="00:05:07.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.76" />
                    <SPLIT distance="100" swimtime="00:02:25.20" />
                    <SPLIT distance="150" swimtime="00:03:42.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="380" reactiontime="+109" swimtime="00:08:01.14" resultid="41747" heatid="45009" lane="6" entrytime="00:07:51.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.83" />
                    <SPLIT distance="100" swimtime="00:01:53.30" />
                    <SPLIT distance="150" swimtime="00:02:56.89" />
                    <SPLIT distance="200" swimtime="00:03:58.66" />
                    <SPLIT distance="250" swimtime="00:05:00.56" />
                    <SPLIT distance="300" swimtime="00:06:01.53" />
                    <SPLIT distance="350" swimtime="00:07:04.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Goncalo Jorge" lastname="Caldeira" birthdate="1996-01-11" gender="M" nation="POR" license="214023" swrid="5464032" athleteid="41730">
              <RESULTS>
                <RESULT eventid="1058" points="375" swimtime="00:12:02.36" resultid="41731" heatid="45085" lane="7" entrytime="00:11:02.92">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.06" />
                    <SPLIT distance="200" swimtime="00:02:45.78" />
                    <SPLIT distance="300" swimtime="00:04:18.36" />
                    <SPLIT distance="400" swimtime="00:05:52.14" />
                    <SPLIT distance="500" swimtime="00:07:25.38" />
                    <SPLIT distance="600" swimtime="00:09:00.62" />
                    <SPLIT distance="700" swimtime="00:10:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="536" reactiontime="+74" swimtime="00:00:30.85" resultid="41732" heatid="44898" lane="3" entrytime="00:00:31.36" />
                <RESULT eventid="2323" points="452" reactiontime="+72" swimtime="00:01:14.07" resultid="41733" heatid="44928" lane="3" entrytime="00:01:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="474" reactiontime="+82" swimtime="00:01:06.31" resultid="41734" heatid="45112" lane="5" entrytime="00:01:05.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="369" reactiontime="+71" swimtime="00:05:49.75" resultid="41735" heatid="45130" lane="5" entrytime="00:05:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                    <SPLIT distance="100" swimtime="00:01:15.13" />
                    <SPLIT distance="150" swimtime="00:01:59.39" />
                    <SPLIT distance="200" swimtime="00:02:44.81" />
                    <SPLIT distance="250" swimtime="00:03:33.39" />
                    <SPLIT distance="300" swimtime="00:04:19.72" />
                    <SPLIT distance="350" swimtime="00:05:05.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="LAGAC" nation="POR" region="ANALG" clubid="41932" swrid="81585" name="Lagoa Academico Clube" shortname="Lagoa AC">
          <ATHLETES>
            <ATHLETE firstname="Filipe Bjorcke" lastname="Santos" birthdate="1988-06-08" gender="M" nation="POR" license="123823" swrid="4781258" athleteid="41948">
              <HANDICAP breast="21" free="21" medley="21" />
              <RESULTS>
                <RESULT eventid="2682" points="398" reactiontime="+81" swimtime="00:00:33.99" resultid="41949" heatid="44896" lane="4" entrytime="00:00:35.30" entrycourse="LCM" />
                <RESULT eventid="2323" points="306" reactiontime="+83" swimtime="00:01:24.12" resultid="41950" heatid="44927" lane="1" entrytime="00:01:22.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="281" reactiontime="+83" swimtime="00:01:17.56" resultid="41951" heatid="45108" lane="6" entrytime="00:01:18.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="210" reactiontime="+105" swimtime="00:00:43.77" resultid="41952" heatid="45018" lane="5" entrytime="00:00:41.18" entrycourse="LCM" />
                <RESULT eventid="2652" points="359" reactiontime="+85" swimtime="00:00:32.71" resultid="41953" heatid="45040" lane="8" entrytime="00:00:32.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Bernardo" lastname="Barbara" birthdate="1970-04-20" gender="F" nation="POR" license="116656" swrid="4432493" athleteid="41933">
              <RESULTS>
                <RESULT eventid="1060" points="250" swimtime="00:15:39.61" resultid="41934" heatid="45075" lane="5" entrytime="00:15:57.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.50" />
                    <SPLIT distance="200" swimtime="00:03:39.67" />
                    <SPLIT distance="300" swimtime="00:05:43.08" />
                    <SPLIT distance="400" swimtime="00:07:46.82" />
                    <SPLIT distance="500" swimtime="00:09:48.18" />
                    <SPLIT distance="600" swimtime="00:11:48.47" />
                    <SPLIT distance="700" swimtime="00:13:46.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2203" points="332" reactiontime="+78" swimtime="00:01:48.89" resultid="41935" heatid="44881" lane="1" entrytime="00:02:00.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2308" points="360" reactiontime="+71" swimtime="00:03:50.50" resultid="41936" heatid="44914" lane="8" entrytime="00:04:06.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.39" />
                    <SPLIT distance="100" swimtime="00:01:53.01" />
                    <SPLIT distance="150" swimtime="00:02:54.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2552" points="251" reactiontime="+90" swimtime="00:01:53.13" resultid="41937" heatid="44922" lane="6" entrytime="00:02:14.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="268" reactiontime="+88" swimtime="00:07:27.02" resultid="41938" heatid="45009" lane="2" entrytime="00:07:52.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.37" />
                    <SPLIT distance="100" swimtime="00:01:42.03" />
                    <SPLIT distance="150" swimtime="00:02:39.80" />
                    <SPLIT distance="200" swimtime="00:03:39.13" />
                    <SPLIT distance="250" swimtime="00:04:38.21" />
                    <SPLIT distance="300" swimtime="00:05:36.78" />
                    <SPLIT distance="350" swimtime="00:06:32.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena Isabel" lastname="Ribeiro" birthdate="1974-02-15" gender="F" nation="POR" license="122493" swrid="4721191" athleteid="41943">
              <RESULTS>
                <RESULT eventid="1060" points="229" swimtime="00:15:48.08" resultid="41944" heatid="45076" lane="7" entrytime="00:15:30.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.60" />
                    <SPLIT distance="200" swimtime="00:03:47.94" />
                    <SPLIT distance="300" swimtime="00:05:47.91" />
                    <SPLIT distance="400" swimtime="00:07:49.45" />
                    <SPLIT distance="500" swimtime="00:09:49.91" />
                    <SPLIT distance="600" swimtime="00:11:51.14" />
                    <SPLIT distance="700" swimtime="00:13:51.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="295" reactiontime="+75" swimtime="00:01:30.00" resultid="41945" heatid="44955" lane="8" entrytime="00:01:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="247" reactiontime="+83" swimtime="00:07:32.89" resultid="41946" heatid="45010" lane="8" entrytime="00:07:27.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.85" />
                    <SPLIT distance="100" swimtime="00:01:41.94" />
                    <SPLIT distance="150" swimtime="00:02:39.47" />
                    <SPLIT distance="200" swimtime="00:03:37.53" />
                    <SPLIT distance="250" swimtime="00:04:36.09" />
                    <SPLIT distance="300" swimtime="00:05:35.28" />
                    <SPLIT distance="350" swimtime="00:06:35.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="348" reactiontime="+80" swimtime="00:00:39.48" resultid="41947" heatid="45068" lane="3" entrytime="00:00:39.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina Monica" lastname="Silva" birthdate="1967-09-24" gender="F" nation="POR" license="205154" swrid="5231630" athleteid="41959">
              <RESULTS>
                <RESULT eventid="1060" status="WDR" swimtime="00:00:00.00" resultid="41960" entrytime="00:18:12.21" entrycourse="LCM" />
                <RESULT eventid="2173" status="WDR" swimtime="00:00:00.00" resultid="41961" entrytime="00:04:54.58" entrycourse="LCM" />
                <RESULT eventid="2607" status="WDR" swimtime="00:00:00.00" resultid="41962" entrytime="00:00:59.11" entrycourse="LCM" />
                <RESULT eventid="2460" status="WDR" swimtime="00:00:00.00" resultid="41963" entrytime="00:02:17.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Pedro" lastname="Sequeira" birthdate="1977-07-18" gender="M" nation="POR" license="213800" swrid="5456928" athleteid="41954">
              <RESULTS>
                <RESULT eventid="1058" status="WDR" swimtime="00:00:00.00" resultid="41955" entrytime="00:15:45.00" />
                <RESULT eventid="2507" status="WDR" swimtime="00:00:00.00" resultid="41956" entrytime="00:03:50.00" />
                <RESULT eventid="2415" status="WDR" swimtime="00:00:00.00" resultid="41957" entrytime="00:01:50.00" />
                <RESULT eventid="2263" status="WDR" swimtime="00:00:00.00" resultid="41958" entrytime="00:07:40.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcia Silva" lastname="Nunes" birthdate="1975-09-14" gender="F" nation="POR" license="122495" swrid="4721190" athleteid="41939">
              <RESULTS>
                <RESULT eventid="2278" status="WDR" swimtime="00:00:00.00" resultid="41940" entrytime="00:04:00.00" />
                <RESULT eventid="2637" status="WDR" swimtime="00:00:00.00" resultid="41941" entrytime="00:01:47.40" />
                <RESULT eventid="2430" status="WDR" swimtime="00:00:00.00" resultid="41942" entrytime="00:00:44.94" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo Alexandre" lastname="Sousa" birthdate="1972-05-16" gender="M" nation="POR" license="106650" swrid="4313167" athleteid="41964">
              <RESULTS>
                <RESULT eventid="1058" points="440" swimtime="00:11:36.64" resultid="41965" heatid="45084" lane="4" entrytime="00:11:09.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.96" />
                    <SPLIT distance="200" swimtime="00:02:44.94" />
                    <SPLIT distance="300" swimtime="00:04:12.34" />
                    <SPLIT distance="400" swimtime="00:05:41.00" />
                    <SPLIT distance="500" swimtime="00:07:10.23" />
                    <SPLIT distance="600" swimtime="00:08:40.60" />
                    <SPLIT distance="700" swimtime="00:10:10.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="464" reactiontime="+94" swimtime="00:02:34.09" resultid="41966" heatid="45094" lane="7" entrytime="00:02:31.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                    <SPLIT distance="100" swimtime="00:01:13.57" />
                    <SPLIT distance="150" swimtime="00:01:52.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="437" reactiontime="+98" swimtime="00:03:01.38" resultid="41967" heatid="44978" lane="7" entrytime="00:03:10.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                    <SPLIT distance="100" swimtime="00:01:21.78" />
                    <SPLIT distance="150" swimtime="00:02:16.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="461" reactiontime="+114" swimtime="00:05:31.47" resultid="41968" heatid="45130" lane="6" entrytime="00:05:22.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                    <SPLIT distance="100" swimtime="00:01:17.42" />
                    <SPLIT distance="150" swimtime="00:01:59.39" />
                    <SPLIT distance="200" swimtime="00:02:41.44" />
                    <SPLIT distance="250" swimtime="00:03:24.39" />
                    <SPLIT distance="300" swimtime="00:04:07.42" />
                    <SPLIT distance="350" swimtime="00:04:50.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="454" reactiontime="+113" swimtime="00:06:33.20" resultid="41969" heatid="45061" lane="7" entrytime="00:06:27.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                    <SPLIT distance="100" swimtime="00:01:31.59" />
                    <SPLIT distance="150" swimtime="00:02:25.00" />
                    <SPLIT distance="200" swimtime="00:03:18.02" />
                    <SPLIT distance="250" swimtime="00:04:17.18" />
                    <SPLIT distance="300" swimtime="00:05:13.62" />
                    <SPLIT distance="350" swimtime="00:05:54.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Susana Matias" lastname="Trindade" birthdate="1974-03-06" gender="F" nation="POR" license="141445" swrid="5125102" athleteid="41970">
              <RESULTS>
                <RESULT eventid="2338" points="427" reactiontime="+86" swimtime="00:00:40.04" resultid="41971" heatid="44890" lane="4" entrytime="00:00:40.42" entrycourse="LCM" />
                <RESULT eventid="2637" points="411" reactiontime="+90" swimtime="00:01:20.58" resultid="41972" heatid="44954" lane="4" entrytime="00:01:29.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="538" reactiontime="+90" swimtime="00:00:34.14" resultid="41973" heatid="45070" lane="6" entrytime="00:00:35.50" entrycourse="LCM" />
                <RESULT eventid="2203" points="341" reactiontime="+75" swimtime="00:01:40.73" resultid="41974" heatid="44883" lane="8" entrytime="00:01:30.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CAPGE" nation="POR" region="ANCNP" clubid="42440" swrid="65876" name="Assoc Pais Amigos Criancas Gaf da Encarnacao" shortname="Gafanha da Encarnacao">
          <ATHLETES>
            <ATHLETE firstname="Rodrigo Alexandre" lastname="Ramos" birthdate="1986-04-24" gender="M" nation="BRA" license="210469" swrid="5361370" athleteid="42447">
              <RESULTS>
                <RESULT eventid="2188" points="192" reactiontime="+100" swimtime="00:00:50.63" resultid="42448" heatid="44941" lane="2" entrytime="00:00:48.83" />
                <RESULT eventid="2415" points="260" reactiontime="+88" swimtime="00:01:21.41" resultid="42449" heatid="45108" lane="1" entrytime="00:01:20.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="194" reactiontime="+90" swimtime="00:01:54.74" resultid="42450" heatid="44994" lane="1" entrytime="00:01:44.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana Cabral" lastname="Oliveira" birthdate="1985-06-30" gender="F" nation="POR" license="131965" swrid="5045154" athleteid="42444">
              <RESULTS>
                <RESULT eventid="2492" status="DNS" swimtime="00:00:00.00" resultid="42445" heatid="45012" lane="7" entrytime="00:06:23.72" />
                <RESULT eventid="2430" status="DNS" swimtime="00:00:00.00" resultid="42446" heatid="45069" lane="6" entrytime="00:00:38.24" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Manuela" lastname="Sequeira" birthdate="1968-08-13" gender="F" nation="POR" license="109962" swrid="4372593" athleteid="42457">
              <RESULTS>
                <RESULT eventid="2308" points="436" reactiontime="+100" swimtime="00:03:36.28" resultid="42458" heatid="44914" lane="3" entrytime="00:03:37.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.03" />
                    <SPLIT distance="100" swimtime="00:01:46.27" />
                    <SPLIT distance="150" swimtime="00:02:42.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2607" points="587" reactiontime="+91" swimtime="00:00:43.84" resultid="42459" heatid="45102" lane="2" entrytime="00:00:43.70" entrycourse="LCM" />
                <RESULT eventid="2460" points="606" reactiontime="+93" swimtime="00:01:38.08" resultid="42460" heatid="45122" lane="5" entrytime="00:01:37.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara Rocha" lastname="Vieira" birthdate="1994-08-17" gender="F" nation="POR" license="207020" swrid="5344269" athleteid="42461">
              <RESULTS>
                <RESULT eventid="1060" points="288" swimtime="00:13:56.32" resultid="42462" heatid="45077" lane="4" entrytime="00:13:00.01">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.34" />
                    <SPLIT distance="200" swimtime="00:03:21.05" />
                    <SPLIT distance="300" swimtime="00:05:07.71" />
                    <SPLIT distance="400" swimtime="00:06:55.44" />
                    <SPLIT distance="500" swimtime="00:08:44.06" />
                    <SPLIT distance="600" swimtime="00:10:30.37" />
                    <SPLIT distance="700" swimtime="00:12:15.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2278" points="329" reactiontime="+83" swimtime="00:03:05.03" resultid="42463" heatid="44903" lane="4" entrytime="00:03:09.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.58" />
                    <SPLIT distance="100" swimtime="00:01:29.43" />
                    <SPLIT distance="150" swimtime="00:02:17.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="325" reactiontime="+86" swimtime="00:01:23.22" resultid="42464" heatid="44955" lane="2" entrytime="00:01:26.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="316" reactiontime="+88" swimtime="00:06:36.16" resultid="42465" heatid="45011" lane="5" entrytime="00:06:34.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.78" />
                    <SPLIT distance="100" swimtime="00:01:33.62" />
                    <SPLIT distance="150" swimtime="00:02:25.15" />
                    <SPLIT distance="200" swimtime="00:03:16.06" />
                    <SPLIT distance="250" swimtime="00:04:06.92" />
                    <SPLIT distance="300" swimtime="00:04:57.48" />
                    <SPLIT distance="350" swimtime="00:05:47.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Rita" lastname="Ribau" birthdate="1995-06-17" gender="F" nation="POR" license="102808" swrid="4229162" athleteid="42451">
              <RESULTS>
                <RESULT eventid="2203" points="626" reactiontime="+70" swimtime="00:01:17.70" resultid="42452" heatid="44883" lane="6" entrytime="00:01:18.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2278" points="688" reactiontime="+81" swimtime="00:02:24.65" resultid="42453" heatid="44905" lane="3" entrytime="00:02:24.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                    <SPLIT distance="100" swimtime="00:01:09.78" />
                    <SPLIT distance="150" swimtime="00:01:47.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2637" points="668" reactiontime="+82" swimtime="00:01:05.48" resultid="42454" heatid="44955" lane="5" entrytime="00:01:20.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="659" reactiontime="+82" swimtime="00:05:10.08" resultid="42455" heatid="45013" lane="2" entrytime="00:05:32.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                    <SPLIT distance="100" swimtime="00:01:13.00" />
                    <SPLIT distance="150" swimtime="00:01:51.71" />
                    <SPLIT distance="200" swimtime="00:02:31.59" />
                    <SPLIT distance="250" swimtime="00:03:11.41" />
                    <SPLIT distance="300" swimtime="00:03:51.71" />
                    <SPLIT distance="350" swimtime="00:04:31.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="628" reactiontime="+79" swimtime="00:00:30.47" resultid="42456" heatid="45072" lane="6" entrytime="00:00:31.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina Ferreira" lastname="Matos" birthdate="1991-06-20" gender="F" nation="POR" license="203814" swrid="4133125" athleteid="42441">
              <RESULTS>
                <RESULT eventid="2308" points="413" reactiontime="+97" swimtime="00:03:12.61" resultid="42442" heatid="44915" lane="1" entrytime="00:03:12.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.59" />
                    <SPLIT distance="100" swimtime="00:01:35.55" />
                    <SPLIT distance="150" swimtime="00:02:24.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2233" points="416" reactiontime="+97" swimtime="00:03:12.73" resultid="42443" heatid="44973" lane="7" entrytime="00:03:14.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                    <SPLIT distance="100" swimtime="00:01:31.11" />
                    <SPLIT distance="150" swimtime="00:02:27.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CFV" nation="POR" region="ANNP" clubid="42761" swrid="65889" name="Clube Fluvial Vilacondense" shortname="Vilacondense">
          <ATHLETES>
            <ATHLETE firstname="Bruno Santos" lastname="Maia" birthdate="1981-08-09" gender="M" nation="POR" license="212423" swrid="5424166" athleteid="42762">
              <RESULTS>
                <RESULT eventid="2682" points="513" reactiontime="+81" swimtime="00:00:32.35" resultid="42763" heatid="44898" lane="7" entrytime="00:00:31.81" />
                <RESULT eventid="2263" points="560" reactiontime="+89" swimtime="00:05:08.52" resultid="42764" heatid="45130" lane="2" entrytime="00:05:25.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                    <SPLIT distance="100" swimtime="00:01:12.30" />
                    <SPLIT distance="150" swimtime="00:01:50.04" />
                    <SPLIT distance="200" swimtime="00:02:28.81" />
                    <SPLIT distance="250" swimtime="00:03:07.80" />
                    <SPLIT distance="300" swimtime="00:03:48.22" />
                    <SPLIT distance="350" swimtime="00:04:28.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Miguel" lastname="Neves" birthdate="1985-09-28" gender="M" nation="POR" license="23046" swrid="4064361" athleteid="42765">
              <RESULTS>
                <RESULT eventid="2323" points="620" reactiontime="+78" swimtime="00:01:08.28" resultid="42766" heatid="44927" lane="4" entrytime="00:01:18.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="485" reactiontime="+81" swimtime="00:01:06.14" resultid="42767" heatid="45111" lane="1" entrytime="00:01:09.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2567" status="RJC" swimtime="00:00:00.00" resultid="42768" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="INDANC" nation="POR" region="ANC" clubid="42504" swrid="76778" name="Individual ANC">
          <ATHLETES>
            <ATHLETE firstname="Joana Margarida" lastname="Cavaleiro" birthdate="1978-04-29" gender="F" nation="POR" license="209719" swrid="5344176" athleteid="42505">
              <RESULTS>
                <RESULT eventid="2607" points="440" reactiontime="+89" swimtime="00:00:45.96" resultid="42506" heatid="45101" lane="4" entrytime="00:00:44.37" entrycourse="LCM" />
                <RESULT eventid="2637" points="376" reactiontime="+83" swimtime="00:01:23.56" resultid="42507" heatid="44955" lane="6" entrytime="00:01:25.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2492" points="398" reactiontime="+89" swimtime="00:06:24.13" resultid="42508" heatid="45011" lane="3" entrytime="00:06:48.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:29.46" />
                    <SPLIT distance="150" swimtime="00:02:18.39" />
                    <SPLIT distance="200" swimtime="00:03:07.90" />
                    <SPLIT distance="250" swimtime="00:03:57.46" />
                    <SPLIT distance="300" swimtime="00:04:47.20" />
                    <SPLIT distance="350" swimtime="00:05:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="451" reactiontime="+88" swimtime="00:01:40.13" resultid="42509" heatid="45122" lane="1" entrytime="00:01:38.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="417" reactiontime="+87" swimtime="00:00:36.73" resultid="42510" heatid="45069" lane="5" entrytime="00:00:36.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CNPO" nation="POR" region="ANNP" clubid="41616" swrid="73271" name="Clube Naval Povoense" shortname="Naval Povoense">
          <ATHLETES>
            <ATHLETE firstname="Maria Rosa" lastname="Serra" birthdate="1977-05-27" gender="F" nation="POR" license="205535" swrid="5260600" athleteid="41620">
              <RESULTS>
                <RESULT eventid="2607" points="227" reactiontime="+96" swimtime="00:00:57.27" resultid="41621" heatid="45098" lane="2" entrytime="00:00:59.44" />
                <RESULT eventid="2637" points="150" reactiontime="+98" swimtime="00:01:53.37" resultid="41622" heatid="44952" lane="3" entrytime="00:01:57.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2460" points="220" reactiontime="+113" swimtime="00:02:07.13" resultid="41623" heatid="45118" lane="4" entrytime="00:02:06.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2430" points="207" reactiontime="+105" swimtime="00:00:46.36" resultid="41624" heatid="45067" lane="2" entrytime="00:00:45.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="David Pereyra" lastname="Noya" birthdate="1975-08-08" gender="M" nation="BOL" license="213527" swrid="5450745" athleteid="41617">
              <RESULTS>
                <RESULT eventid="2188" status="DNS" swimtime="00:00:00.00" resultid="41618" heatid="44939" lane="1" entrytime="00:01:00.00" />
                <RESULT eventid="2293" status="DNS" swimtime="00:00:00.00" resultid="41619" heatid="45015" lane="4" entrytime="00:00:55.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marco Paulo" lastname="Silva" birthdate="1970-10-20" gender="M" nation="POR" license="118005" swrid="4577120" athleteid="41625">
              <RESULTS>
                <RESULT eventid="2622" points="366" reactiontime="+94" swimtime="00:03:43.70" resultid="41626" heatid="44875" lane="8" entrytime="00:03:47.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.99" />
                    <SPLIT distance="100" swimtime="00:01:44.77" />
                    <SPLIT distance="150" swimtime="00:02:45.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="406" reactiontime="+97" swimtime="00:01:16.78" resultid="41627" heatid="45108" lane="2" entrytime="00:01:18.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="357" reactiontime="+100" swimtime="00:01:42.11" resultid="41628" heatid="44994" lane="5" entrytime="00:01:42.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="374" reactiontime="+87" swimtime="00:00:43.18" resultid="41629" heatid="44945" lane="7" entrytime="00:00:42.79" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="VNC" nation="POR" region="ANMIN" clubid="43574" swrid="65810" name="Viana Natacao Clube" shortname="Viana Natacao">
          <ATHLETES>
            <ATHLETE firstname="Rui Miguel" lastname="Pinto" birthdate="1969-03-22" gender="M" nation="POR" license="106906" swrid="5115794" athleteid="43589">
              <RESULTS>
                <RESULT eventid="2507" status="DNS" swimtime="00:00:00.00" resultid="43590" heatid="45091" lane="6" entrytime="00:03:23.19" entrycourse="LCM" />
                <RESULT eventid="2188" points="339" reactiontime="+102" swimtime="00:00:44.61" resultid="43591" heatid="44942" lane="4" entrytime="00:00:45.42" entrycourse="LCM" />
                <RESULT eventid="2415" points="340" reactiontime="+100" swimtime="00:01:21.40" resultid="43592" heatid="45107" lane="4" entrytime="00:01:21.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="377" reactiontime="+101" swimtime="00:00:34.75" resultid="43593" heatid="45038" lane="5" entrytime="00:00:33.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos Alberto" lastname="Couteiro" birthdate="1945-10-20" gender="M" nation="POR" license="201514" swrid="5171428" athleteid="43579">
              <RESULTS>
                <RESULT eventid="2537" points="141" reactiontime="+75" swimtime="00:02:38.44" resultid="43580" heatid="44884" lane="6" entrytime="00:02:30.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:13.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2218" points="136" reactiontime="+101" swimtime="00:05:48.74" resultid="43581" heatid="44916" lane="3" entrytime="00:05:45.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.84" />
                    <SPLIT distance="100" swimtime="00:02:46.31" />
                    <SPLIT distance="150" swimtime="00:04:18.65" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="716 - Durante o percurso não rodou os pés para fora durante a parte propulsiva da pernada - SW 7.5" eventid="2445" reactiontime="+135" status="DSQ" swimtime="00:02:26.57" resultid="43582" heatid="44990" lane="6" entrytime="00:02:26.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="181" reactiontime="+81" swimtime="00:01:05.72" resultid="43583" heatid="45014" lane="7" entrytime="00:01:10.50" />
                <RESULT eventid="2652" points="161" reactiontime="+118" swimtime="00:00:57.32" resultid="43584" heatid="45032" lane="5" entrytime="00:01:05.50" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ivone Dorinda" lastname="Silva" birthdate="1975-03-14" gender="F" nation="POR" license="14420" swrid="4575823" athleteid="43594">
              <RESULTS>
                <RESULT eventid="2522" status="DNS" swimtime="00:00:00.00" resultid="43595" heatid="45026" lane="4" entrytime="00:00:38.57" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Eduardo" lastname="Couteiro" birthdate="1976-05-11" gender="M" nation="POR" license="106905" swrid="5032034" athleteid="43585">
              <RESULTS>
                <RESULT eventid="2682" points="778" reactiontime="+77" swimtime="00:00:28.87" resultid="43586" heatid="44898" lane="1" entrytime="00:00:31.92" entrycourse="LCM" />
                <RESULT eventid="2188" points="739" reactiontime="+74" swimtime="00:00:33.07" resultid="43587" heatid="44949" lane="4" entrytime="00:00:35.09" entrycourse="LCM" />
                <RESULT eventid="2293" points="649" reactiontime="+65" swimtime="00:00:33.23" resultid="43588" heatid="45020" lane="2" entrytime="00:00:34.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor Borges" lastname="Carvalho" birthdate="1964-06-14" gender="M" nation="POR" license="14392" swrid="4574566" athleteid="43575">
              <RESULTS>
                <RESULT eventid="2188" points="318" reactiontime="+104" swimtime="00:00:45.46" resultid="43576" heatid="44944" lane="2" entrytime="00:00:44.15" entrycourse="LCM" />
                <RESULT eventid="2415" status="DNS" swimtime="00:00:00.00" resultid="43577" heatid="45108" lane="5" entrytime="00:01:18.25" entrycourse="LCM" />
                <RESULT eventid="2445" status="DNS" swimtime="00:00:00.00" resultid="43578" heatid="44993" lane="6" entrytime="00:01:47.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SAD" nation="POR" region="ANL" clubid="41650" swrid="65806" name="Sport Alges e Dafundo" shortname="Alges">
          <ATHLETES>
            <ATHLETE firstname="Jose Manuel" lastname="Horta" birthdate="1949-08-21" gender="M" nation="POR" license="141654" swrid="5119298" athleteid="41675">
              <RESULTS>
                <RESULT eventid="2622" points="187" swimtime="00:05:36.53" resultid="41676" heatid="44872" lane="3" entrytime="00:05:29.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.27" />
                    <SPLIT distance="100" swimtime="00:02:46.67" />
                    <SPLIT distance="150" swimtime="00:04:14.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="198" reactiontime="+119" swimtime="00:01:03.18" resultid="41677" heatid="44938" lane="6" entrytime="00:01:02.98" entrycourse="LCM" />
                <RESULT eventid="2263" points="86" reactiontime="+124" swimtime="00:12:16.04" resultid="41678" heatid="45124" lane="2" entrytime="00:11:08.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.11" />
                    <SPLIT distance="100" swimtime="00:02:48.77" />
                    <SPLIT distance="150" swimtime="00:04:25.11" />
                    <SPLIT distance="200" swimtime="00:06:03.05" />
                    <SPLIT distance="250" swimtime="00:07:37.16" />
                    <SPLIT distance="300" swimtime="00:09:12.91" />
                    <SPLIT distance="350" swimtime="00:10:45.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2445" points="164" reactiontime="+129" swimtime="00:02:36.51" resultid="41679" heatid="44990" lane="2" entrytime="00:02:28.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="101" reactiontime="+122" swimtime="00:01:00.99" resultid="41680" heatid="45033" lane="6" entrytime="00:00:54.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos Manuel" lastname="Lopes" birthdate="1966-03-05" gender="M" nation="POR" license="202483" swrid="4797614" athleteid="41669">
              <RESULTS>
                <RESULT eventid="2218" points="100" reactiontime="+92" swimtime="00:05:24.61" resultid="41670" heatid="44916" lane="5" entrytime="00:05:27.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.94" />
                    <SPLIT distance="100" swimtime="00:02:34.55" />
                    <SPLIT distance="150" swimtime="00:04:03.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2323" points="96" reactiontime="+95" swimtime="00:02:20.85" resultid="41671" heatid="44925" lane="6" entrytime="00:02:11.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="159" reactiontime="+92" swimtime="00:04:42.28" resultid="41672" heatid="44975" lane="6" entrytime="00:04:40.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.40" />
                    <SPLIT distance="100" swimtime="00:02:21.08" />
                    <SPLIT distance="150" swimtime="00:03:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="823 - efectuou duas pernadas por cada ciclo de braçada - MSW 3.9" eventid="2567" reactiontime="+89" status="DSQ" swimtime="00:05:37.42" resultid="41673" heatid="45028" lane="3" entrytime="00:04:58.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.53" />
                    <SPLIT distance="100" swimtime="00:02:25.86" />
                    <SPLIT distance="150" swimtime="00:03:55.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2248" points="147" reactiontime="+94" swimtime="00:10:26.05" resultid="41674" heatid="45058" lane="3" entrytime="00:10:35.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.23" />
                    <SPLIT distance="100" swimtime="00:02:19.86" />
                    <SPLIT distance="150" swimtime="00:03:52.33" />
                    <SPLIT distance="200" swimtime="00:05:18.17" />
                    <SPLIT distance="250" swimtime="00:06:40.25" />
                    <SPLIT distance="300" swimtime="00:08:03.77" />
                    <SPLIT distance="350" swimtime="00:09:14.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Maria" lastname="Ferreira" birthdate="1950-07-20" gender="F" nation="POR" license="100434" swrid="4224012" athleteid="41706">
              <RESULTS>
                <RESULT eventid="2522" status="DNS" swimtime="00:00:00.00" resultid="41707" heatid="45024" lane="3" entrytime="00:00:51.02" entrycourse="LCM" />
                <RESULT eventid="2430" status="DNS" swimtime="00:00:00.00" resultid="41708" heatid="45068" lane="4" entrytime="00:00:39.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Vidigal" lastname="Salgueiro" birthdate="1945-07-07" gender="M" nation="POR" license="119671" swrid="4610259" athleteid="41651">
              <RESULTS>
                <RESULT eventid="1058" status="DNF" swimtime="00:00:00.00" resultid="41652" heatid="45080" lane="6" entrytime="00:16:53.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:03.46" />
                    <SPLIT distance="200" swimtime="00:04:16.52" />
                    <SPLIT distance="300" swimtime="00:06:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="356" swimtime="00:03:45.51" resultid="41653" heatid="45090" lane="4" entrytime="00:03:39.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.36" />
                    <SPLIT distance="100" swimtime="00:01:48.35" />
                    <SPLIT distance="150" swimtime="00:02:51.74" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rec Nac Esc K" eventid="2415" points="436" swimtime="00:01:34.65" resultid="41654" heatid="45105" lane="7" entrytime="00:01:33.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="307" swimtime="00:08:29.67" resultid="41655" heatid="45125" lane="6" entrytime="00:07:55.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.85" />
                    <SPLIT distance="100" swimtime="00:02:05.32" />
                    <SPLIT distance="150" swimtime="00:03:13.30" />
                    <SPLIT distance="200" swimtime="00:04:19.07" />
                    <SPLIT distance="250" swimtime="00:05:25.97" />
                    <SPLIT distance="300" swimtime="00:06:30.50" />
                    <SPLIT distance="350" swimtime="00:07:34.50" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rec Nac Esc K" eventid="2652" points="461" reactiontime="+117" swimtime="00:00:40.37" resultid="41656" heatid="45035" lane="3" entrytime="00:00:39.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jaime Carlos" lastname="Bento" birthdate="1961-03-05" gender="M" nation="POR" license="118614" swrid="4583590" athleteid="41683">
              <RESULTS>
                <RESULT comment="Rec Nac Esc H" eventid="1058" points="832" swimtime="00:11:05.20" resultid="41684" heatid="45084" lane="6" entrytime="00:11:30.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.06" />
                    <SPLIT distance="200" swimtime="00:02:42.20" />
                    <SPLIT distance="300" swimtime="00:04:06.21" />
                    <SPLIT distance="400" swimtime="00:05:30.66" />
                    <SPLIT distance="500" swimtime="00:06:55.46" />
                    <SPLIT distance="600" swimtime="00:08:19.62" />
                    <SPLIT distance="700" swimtime="00:09:43.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2507" points="797" reactiontime="+94" swimtime="00:02:30.86" resultid="41685" heatid="45094" lane="2" entrytime="00:02:31.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:13.59" />
                    <SPLIT distance="150" swimtime="00:01:52.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="718" reactiontime="+95" swimtime="00:01:08.15" resultid="41686" heatid="45111" lane="6" entrytime="00:01:08.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="766" reactiontime="+96" swimtime="00:05:27.62" resultid="41687" heatid="45130" lane="1" entrytime="00:05:33.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:15.03" />
                    <SPLIT distance="150" swimtime="00:01:55.50" />
                    <SPLIT distance="200" swimtime="00:02:38.11" />
                    <SPLIT distance="250" swimtime="00:03:20.88" />
                    <SPLIT distance="300" swimtime="00:04:03.75" />
                    <SPLIT distance="350" swimtime="00:04:46.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="695" reactiontime="+92" swimtime="00:00:30.85" resultid="41688" heatid="45041" lane="4" entrytime="00:00:30.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Manuel" lastname="Ferreira" birthdate="1948-11-19" gender="M" nation="POR" license="123326" swrid="4756577" athleteid="41712">
              <RESULTS>
                <RESULT eventid="2293" status="DNS" swimtime="00:00:00.00" resultid="41713" heatid="45014" lane="3" entrytime="00:01:05.02" entrycourse="LCM" />
                <RESULT eventid="2652" status="DNS" swimtime="00:00:00.00" resultid="41714" heatid="45032" lane="3" entrytime="00:01:10.21" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor Manuel" lastname="Mavioso" birthdate="1956-11-11" gender="M" nation="POR" license="100689" swrid="4800291" athleteid="41692">
              <RESULTS>
                <RESULT comment="Rec Nac Esc I" eventid="2218" points="674" reactiontime="+86" swimtime="00:03:03.56" resultid="41693" heatid="44920" lane="7" entrytime="00:03:00.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.80" />
                    <SPLIT distance="100" swimtime="00:01:29.51" />
                    <SPLIT distance="150" swimtime="00:02:17.97" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rec Nac Esc I" eventid="2323" points="733" reactiontime="+98" swimtime="00:01:21.08" resultid="41694" heatid="44927" lane="3" entrytime="00:01:20.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="465" reactiontime="+80" swimtime="00:00:44.54" resultid="41695" heatid="44941" lane="4" entrytime="00:00:47.23" entrycourse="SCM" />
                <RESULT comment="Rec Nac Esc I" eventid="2415" points="770" reactiontime="+78" swimtime="00:01:08.48" resultid="41696" heatid="45111" lane="7" entrytime="00:01:09.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Rec Nac Esc I" eventid="2385" points="793" reactiontime="+90" swimtime="00:02:58.90" resultid="41697" heatid="44979" lane="5" entrytime="00:02:56.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:22.93" />
                    <SPLIT distance="150" swimtime="00:02:20.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Jose" lastname="Trabuco" birthdate="1950-07-04" gender="M" nation="POR" license="148719" swrid="5106730" athleteid="41681">
              <RESULTS>
                <RESULT eventid="2652" points="576" reactiontime="+95" swimtime="00:00:34.20" resultid="41682" heatid="45039" lane="6" entrytime="00:00:33.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre Azevedo" lastname="Gaspar" birthdate="1945-04-08" gender="M" nation="POR" license="119670" swrid="4610230" athleteid="41663">
              <RESULTS>
                <RESULT comment="Rec Nac Esc K" eventid="2622" points="499" reactiontime="+115" swimtime="00:04:17.23" resultid="41664" heatid="44874" lane="8" entrytime="00:04:18.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.70" />
                    <SPLIT distance="100" swimtime="00:02:04.55" />
                    <SPLIT distance="150" swimtime="00:03:11.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="438" reactiontime="+114" swimtime="00:00:52.08" resultid="41665" heatid="44940" lane="2" entrytime="00:00:51.03" entrycourse="LCM" />
                <RESULT comment="Rec Nac Esc K" eventid="2385" points="335" reactiontime="+121" swimtime="00:04:29.60" resultid="41666" heatid="44975" lane="3" entrytime="00:04:11.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.51" />
                    <SPLIT distance="100" swimtime="00:02:17.57" />
                    <SPLIT distance="150" swimtime="00:03:24.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2293" points="262" reactiontime="+88" swimtime="00:00:58.17" resultid="41667" heatid="45015" lane="1" entrytime="00:00:57.02" entrycourse="LCM" />
                <RESULT eventid="2445" points="417" reactiontime="+100" swimtime="00:02:00.34" resultid="41668" heatid="44992" lane="6" entrytime="00:01:57.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stephen Thomas" lastname="Dyson" birthdate="1947-09-24" gender="M" nation="POR" license="109270" swrid="4345520" athleteid="41657">
              <RESULTS>
                <RESULT eventid="1058" points="696" swimtime="00:13:01.83" resultid="41658" heatid="45082" lane="4" entrytime="00:13:03.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.04" />
                    <SPLIT distance="200" swimtime="00:03:15.23" />
                    <SPLIT distance="300" swimtime="00:04:55.15" />
                    <SPLIT distance="400" swimtime="00:06:33.87" />
                    <SPLIT distance="500" swimtime="00:08:11.51" />
                    <SPLIT distance="600" swimtime="00:09:49.05" />
                    <SPLIT distance="700" swimtime="00:11:26.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2682" points="323" reactiontime="+99" swimtime="00:00:46.02" resultid="41659" heatid="44895" lane="2" entrytime="00:00:39.77" entrycourse="LCM" />
                <RESULT eventid="2507" points="598" reactiontime="+91" swimtime="00:03:01.49" resultid="41660" heatid="45092" lane="5" entrytime="00:02:53.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:25.89" />
                    <SPLIT distance="150" swimtime="00:02:14.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2415" points="557" reactiontime="+99" swimtime="00:01:19.72" resultid="41661" heatid="45108" lane="7" entrytime="00:01:19.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2263" points="653" reactiontime="+100" swimtime="00:06:15.37" resultid="41662" heatid="45128" lane="8" entrytime="00:06:28.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.99" />
                    <SPLIT distance="100" swimtime="00:01:27.22" />
                    <SPLIT distance="150" swimtime="00:02:15.35" />
                    <SPLIT distance="200" swimtime="00:03:03.60" />
                    <SPLIT distance="250" swimtime="00:03:52.36" />
                    <SPLIT distance="300" swimtime="00:04:40.48" />
                    <SPLIT distance="350" swimtime="00:05:28.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo Marcos" lastname="Dantas" birthdate="1963-11-18" gender="M" nation="POR" license="206918" swrid="5276386" athleteid="41715">
              <RESULTS>
                <RESULT eventid="2507" points="595" reactiontime="+71" swimtime="00:02:34.00" resultid="41716" heatid="45094" lane="3" entrytime="00:02:30.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                    <SPLIT distance="100" swimtime="00:01:13.51" />
                    <SPLIT distance="150" swimtime="00:01:53.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="466" reactiontime="+79" swimtime="00:00:40.05" resultid="41717" heatid="44943" lane="1" entrytime="00:00:45.08" />
                <RESULT eventid="2415" points="669" reactiontime="+69" swimtime="00:01:08.70" resultid="41718" heatid="45111" lane="2" entrytime="00:01:09.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2385" points="507" reactiontime="+74" swimtime="00:03:12.07" resultid="41719" heatid="44979" lane="8" entrytime="00:03:05.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                    <SPLIT distance="100" swimtime="00:01:34.50" />
                    <SPLIT distance="150" swimtime="00:02:28.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2652" points="668" reactiontime="+77" swimtime="00:00:30.43" resultid="41720" heatid="45042" lane="6" entrytime="00:00:29.98" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karin" lastname="Potter" birthdate="1959-02-20" gender="F" nation="BRA" license="210165" swrid="5351811" athleteid="41703">
              <RESULTS>
                <RESULT eventid="2522" points="559" reactiontime="+99" swimtime="00:00:47.23" resultid="41704" heatid="45025" lane="8" entrytime="00:00:47.01" entrycourse="LCM" />
                <RESULT comment="810 - Movimento alternado de pernas após viragem aos 50 m - SW 8.3" eventid="2400" status="DSQ" swimtime="00:00:00.00" resultid="41705" heatid="45063" lane="5" entrytime="00:08:30.00" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mario Gomes" lastname="Bairrada" birthdate="1952-08-30" gender="M" nation="POR" license="100885" swrid="4345366" athleteid="41698">
              <RESULTS>
                <RESULT eventid="2622" points="381" reactiontime="+108" swimtime="00:04:18.69" resultid="41699" heatid="44874" lane="3" entrytime="00:03:58.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.26" />
                    <SPLIT distance="100" swimtime="00:02:03.74" />
                    <SPLIT distance="150" swimtime="00:03:11.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2188" points="322" reactiontime="+102" swimtime="00:00:50.32" resultid="41700" heatid="44941" lane="7" entrytime="00:00:49.29" entrycourse="LCM" />
                <RESULT eventid="2385" status="DNS" swimtime="00:00:00.00" resultid="41701" heatid="44976" lane="8" entrytime="00:04:05.07" entrycourse="LCM" />
                <RESULT eventid="2445" status="DNS" swimtime="00:00:00.00" resultid="41702" heatid="44993" lane="7" entrytime="00:01:48.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Felix" lastname="Ferreira" birthdate="1954-01-10" gender="F" nation="POR" license="112081" swrid="4413292" athleteid="41689">
              <RESULTS>
                <RESULT eventid="2607" points="292" reactiontime="+112" swimtime="00:01:02.52" resultid="41690" heatid="45098" lane="8" entrytime="00:01:04.86" entrycourse="LCM" />
                <RESULT eventid="2637" points="176" reactiontime="+106" swimtime="00:02:08.37" resultid="41691" heatid="44952" lane="2" entrytime="00:02:06.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Violante Isabel" lastname="Ribeiro" birthdate="1967-05-11" gender="F" nation="POR" license="124926" swrid="4005228" athleteid="41709">
              <RESULTS>
                <RESULT eventid="2203" status="DNS" swimtime="00:00:00.00" resultid="41710" heatid="44880" lane="4" entrytime="00:02:02.51" entrycourse="LCM" />
                <RESULT eventid="2278" status="DNS" swimtime="00:00:00.00" resultid="41711" heatid="44902" lane="7" entrytime="00:04:31.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
