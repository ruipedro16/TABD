<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Associação de Natação do Norte de Portugal" version="11.71436">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Paços de Ferreira" name="Troféu Pescada - José Carlos Freitas e Troféu Master ANNP" name.en="Troféu Pescada - José Carlos Freitas e Troféu Master ANNP" course="SCM" deadline="2021-11-25" entrystartdate="2021-10-01" entrytype="OPEN" organizer="ANNP " result.url="http://annp.pt/provas2122/07" startmethod="1" timing="AUTOMATIC" type="POR.MNP" withdrawuntil="2021-11-26" nation="POR" maxentriesathlete="3">
      <AGEDATE value="2021-12-04" type="YEAR" />
      <POOL name="Piscina Municipal de Paços de Ferreira " lanemin="1" lanemax="8" />
      <FACILITY city="Paços de Ferreira" name="Piscina Municipal de Paços de Ferreira " nation="POR" />
      <POINTTABLE pointtableid="1124" name="DSV Master Performance Table" version="2020" />
      <CONTACT email="info@annp.pt" name="Rita Fougo" />
      <QUALIFY from="2019-01-01" until="2021-11-29" conversion="FINA_POINTS" />
      <SESSIONS>
        <SESSION date="2021-12-04" daytime="09:00" name="1ª Jornada" number="1" warmupfrom="08:00" warmupuntil="08:45">
          <EVENTS>
            <EVENT eventid="10314" daytime="09:00" gender="X" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="EUR" value="350" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10315" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11848" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10316" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11989" />
                    <RANKING order="2" place="2" resultid="12210" />
                    <RANKING order="3" place="3" resultid="12162" />
                    <RANKING order="4" place="4" resultid="12336" />
                    <RANKING order="5" place="5" resultid="12089" />
                    <RANKING order="6" place="6" resultid="11954" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10317" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12642" />
                    <RANKING order="2" place="2" resultid="11847" />
                    <RANKING order="3" place="3" resultid="12092" />
                    <RANKING order="4" place="4" resultid="12337" />
                    <RANKING order="5" place="5" resultid="12533" />
                    <RANKING order="6" place="6" resultid="12414" />
                    <RANKING order="7" place="-1" resultid="12209" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10318" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12343" />
                    <RANKING order="2" place="2" resultid="11846" />
                    <RANKING order="3" place="3" resultid="12417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10319" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12536" />
                    <RANKING order="2" place="-1" resultid="12347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10320" agemax="319" agemin="280" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="12094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10321" agemax="359" agemin="320" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12727" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12728" daytime="09:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12803" daytime="09:10" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4102" daytime="09:15" gender="F" number="2" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4103" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="4104" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="4105" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="4106" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12057" />
                    <RANKING order="2" place="-1" resultid="11766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4107" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="4108" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="4109" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4110" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="4111" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="4112" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="4113" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="4818" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="4114" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12057" />
                    <RANKING order="2" place="-1" resultid="11766" />
                    <RANKING order="3" place="-1" resultid="11895" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12729" daytime="09:15" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="10455">
                  <FEE currency="EUR" value="400" />
                </TIMESTANDARDREF>
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="4128" daytime="09:45" gender="M" number="3" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4129" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="4130" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11914" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4131" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12673" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4132" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12030" />
                    <RANKING order="2" place="2" resultid="12457" />
                    <RANKING order="3" place="-1" resultid="12062" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4133" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12280" />
                    <RANKING order="2" place="2" resultid="12467" />
                    <RANKING order="3" place="-1" resultid="12042" />
                    <RANKING order="4" place="-1" resultid="11892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4134" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="4135" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12088" />
                    <RANKING order="2" place="2" resultid="12301" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4136" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11898" />
                    <RANKING order="2" place="2" resultid="11887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4137" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4138" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="4139" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="4819" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="4140" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11898" />
                    <RANKING order="2" place="2" resultid="11887" />
                    <RANKING order="3" place="3" resultid="11879" />
                    <RANKING order="4" place="4" resultid="12673" />
                    <RANKING order="5" place="5" resultid="12030" />
                    <RANKING order="6" place="6" resultid="12457" />
                    <RANKING order="7" place="7" resultid="12088" />
                    <RANKING order="8" place="8" resultid="12301" />
                    <RANKING order="9" place="9" resultid="12280" />
                    <RANKING order="10" place="10" resultid="12467" />
                    <RANKING order="11" place="11" resultid="11914" />
                    <RANKING order="12" place="-1" resultid="12042" />
                    <RANKING order="13" place="-1" resultid="12062" />
                    <RANKING order="14" place="-1" resultid="11892" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12730" daytime="09:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12731" daytime="10:15" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="10441">
                  <FEE currency="EUR" value="400" />
                </TIMESTANDARDREF>
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="9605" daytime="10:45" gender="F" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10499" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12631" />
                    <RANKING order="2" place="2" resultid="12647" />
                    <RANKING order="3" place="3" resultid="11816" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10500" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="10501" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12151" />
                    <RANKING order="2" place="2" resultid="11934" />
                    <RANKING order="3" place="-1" resultid="12395" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10502" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12268" />
                    <RANKING order="2" place="2" resultid="11820" />
                    <RANKING order="3" place="3" resultid="11938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10503" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12215" />
                    <RANKING order="2" place="2" resultid="12013" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10504" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12006" />
                    <RANKING order="2" place="2" resultid="12264" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10505" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12521" />
                    <RANKING order="2" place="2" resultid="12297" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10506" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12308" />
                    <RANKING order="2" place="2" resultid="11786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10507" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="10508" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="10509" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10510" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10511" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12631" />
                    <RANKING order="2" place="2" resultid="12647" />
                    <RANKING order="3" place="3" resultid="12215" />
                    <RANKING order="4" place="4" resultid="11816" />
                    <RANKING order="5" place="5" resultid="12268" />
                    <RANKING order="6" place="6" resultid="12013" />
                    <RANKING order="7" place="7" resultid="12521" />
                    <RANKING order="8" place="8" resultid="12297" />
                    <RANKING order="9" place="9" resultid="11820" />
                    <RANKING order="10" place="10" resultid="12151" />
                    <RANKING order="11" place="11" resultid="12006" />
                    <RANKING order="12" place="12" resultid="12308" />
                    <RANKING order="13" place="13" resultid="11938" />
                    <RANKING order="14" place="14" resultid="11786" />
                    <RANKING order="15" place="15" resultid="11934" />
                    <RANKING order="16" place="16" resultid="12264" />
                    <RANKING order="17" place="-1" resultid="12395" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12732" daytime="10:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12733" daytime="10:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12804" daytime="10:55" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="9632" daytime="10:55" gender="M" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10538" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11789" />
                    <RANKING order="2" place="2" resultid="11946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10539" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10540" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="10541" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10542" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12054" />
                    <RANKING order="2" place="2" resultid="12079" />
                    <RANKING order="3" place="3" resultid="11942" />
                    <RANKING order="4" place="-1" resultid="11773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10543" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12220" />
                    <RANKING order="2" place="-1" resultid="12045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10544" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12638" />
                    <RANKING order="2" place="-1" resultid="12289" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10545" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10546" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10547" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="10548" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10549" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10550" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12458" />
                    <RANKING order="2" place="2" resultid="11789" />
                    <RANKING order="3" place="3" resultid="12471" />
                    <RANKING order="4" place="4" resultid="12054" />
                    <RANKING order="5" place="5" resultid="11946" />
                    <RANKING order="6" place="6" resultid="12249" />
                    <RANKING order="7" place="7" resultid="12450" />
                    <RANKING order="8" place="8" resultid="12638" />
                    <RANKING order="9" place="9" resultid="12079" />
                    <RANKING order="10" place="10" resultid="12220" />
                    <RANKING order="11" place="11" resultid="11942" />
                    <RANKING order="12" place="-1" resultid="12289" />
                    <RANKING order="13" place="-1" resultid="11773" />
                    <RANKING order="14" place="-1" resultid="12045" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12734" daytime="10:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12735" daytime="11:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2111" daytime="11:05" gender="F" number="6" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4820" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4821" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="4822" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="4823" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12628" />
                    <RANKING order="2" place="2" resultid="12058" />
                    <RANKING order="3" place="3" resultid="12129" />
                    <RANKING order="4" place="-1" resultid="11767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4824" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4825" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4826" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4827" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="4828" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="4829" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="4830" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="4831" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="4832" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11760" />
                    <RANKING order="2" place="2" resultid="11851" />
                    <RANKING order="3" place="3" resultid="12701" />
                    <RANKING order="4" place="4" resultid="12007" />
                    <RANKING order="5" place="5" resultid="12628" />
                    <RANKING order="6" place="6" resultid="12058" />
                    <RANKING order="7" place="7" resultid="12129" />
                    <RANKING order="8" place="-1" resultid="11767" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12736" daytime="11:05" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2124" daytime="11:10" gender="M" number="7" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4885" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="4886" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="4887" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="12311" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4888" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="4889" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12120" />
                    <RANKING order="2" place="2" resultid="12389" />
                    <RANKING order="3" place="-1" resultid="12080" />
                    <RANKING order="4" place="-1" resultid="12203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4890" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12479" />
                    <RANKING order="2" place="2" resultid="12038" />
                    <RANKING order="3" place="3" resultid="12221" />
                    <RANKING order="4" place="-1" resultid="12035" />
                    <RANKING order="5" place="-1" resultid="12046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4891" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4892" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4893" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="4894" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="4895" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="4896" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="4897" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11899" />
                    <RANKING order="2" place="2" resultid="12479" />
                    <RANKING order="3" place="3" resultid="12038" />
                    <RANKING order="4" place="4" resultid="12120" />
                    <RANKING order="5" place="5" resultid="12389" />
                    <RANKING order="6" place="6" resultid="12221" />
                    <RANKING order="7" place="7" resultid="12514" />
                    <RANKING order="8" place="-1" resultid="12080" />
                    <RANKING order="9" place="-1" resultid="12203" />
                    <RANKING order="10" place="-1" resultid="12035" />
                    <RANKING order="11" place="-1" resultid="12046" />
                    <RANKING order="12" place="-1" resultid="12311" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12737" daytime="11:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12738" daytime="11:15" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="9659" daytime="11:20" gender="F" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10512" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12658" />
                    <RANKING order="2" place="2" resultid="12174" />
                    <RANKING order="3" place="3" resultid="12136" />
                    <RANKING order="4" place="4" resultid="12475" />
                    <RANKING order="5" place="5" resultid="12381" />
                    <RANKING order="6" place="6" resultid="12684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10513" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12190" />
                    <RANKING order="2" place="2" resultid="12188" />
                    <RANKING order="3" place="3" resultid="12315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10514" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12257" />
                    <RANKING order="2" place="2" resultid="12396" />
                    <RANKING order="3" place="3" resultid="12506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10515" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12165" />
                    <RANKING order="2" place="2" resultid="12498" />
                    <RANKING order="3" place="-1" resultid="12578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10516" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="10517" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12404" />
                    <RANKING order="2" place="2" resultid="12143" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10518" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12522" />
                    <RANKING order="2" place="2" resultid="12073" />
                    <RANKING order="3" place="3" resultid="12097" />
                    <RANKING order="4" place="4" resultid="11801" />
                    <RANKING order="5" place="5" resultid="12197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10519" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10520" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="10521" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="12010" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10522" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10523" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10524" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12165" />
                    <RANKING order="2" place="2" resultid="12658" />
                    <RANKING order="3" place="3" resultid="12257" />
                    <RANKING order="4" place="4" resultid="12190" />
                    <RANKING order="5" place="5" resultid="12174" />
                    <RANKING order="6" place="6" resultid="12136" />
                    <RANKING order="7" place="7" resultid="12188" />
                    <RANKING order="8" place="8" resultid="12522" />
                    <RANKING order="9" place="9" resultid="12404" />
                    <RANKING order="10" place="10" resultid="12475" />
                    <RANKING order="11" place="11" resultid="12315" />
                    <RANKING order="12" place="12" resultid="12498" />
                    <RANKING order="13" place="13" resultid="12143" />
                    <RANKING order="14" place="14" resultid="12396" />
                    <RANKING order="15" place="15" resultid="12381" />
                    <RANKING order="16" place="16" resultid="12073" />
                    <RANKING order="17" place="17" resultid="12506" />
                    <RANKING order="18" place="17" resultid="12194" />
                    <RANKING order="19" place="19" resultid="12097" />
                    <RANKING order="20" place="20" resultid="11801" />
                    <RANKING order="21" place="21" resultid="12197" />
                    <RANKING order="22" place="22" resultid="12684" />
                    <RANKING order="23" place="-1" resultid="12010" />
                    <RANKING order="24" place="-1" resultid="12578" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12739" daytime="11:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12740" daytime="11:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12741" daytime="11:25" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="9685" daytime="11:30" gender="M" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="9686" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12654" />
                    <RANKING order="2" place="2" resultid="12369" />
                    <RANKING order="3" place="3" resultid="12231" />
                    <RANKING order="4" place="4" resultid="12359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9687" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12253" />
                    <RANKING order="2" place="2" resultid="11907" />
                    <RANKING order="3" place="3" resultid="12122" />
                    <RANKING order="4" place="4" resultid="12666" />
                    <RANKING order="5" place="5" resultid="12490" />
                    <RANKING order="6" place="-1" resultid="12200" />
                    <RANKING order="7" place="-1" resultid="12420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9688" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12662" />
                    <RANKING order="2" place="2" resultid="12155" />
                    <RANKING order="3" place="3" resultid="12486" />
                    <RANKING order="4" place="4" resultid="12149" />
                    <RANKING order="5" place="-1" resultid="12312" />
                    <RANKING order="6" place="-1" resultid="12607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9689" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11957" />
                    <RANKING order="2" place="2" resultid="12529" />
                    <RANKING order="3" place="3" resultid="12565" />
                    <RANKING order="4" place="4" resultid="12604" />
                    <RANKING order="5" place="5" resultid="12611" />
                    <RANKING order="6" place="6" resultid="12582" />
                    <RANKING order="7" place="7" resultid="11827" />
                    <RANKING order="8" place="8" resultid="12619" />
                    <RANKING order="9" place="-1" resultid="12377" />
                    <RANKING order="10" place="-1" resultid="12401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9690" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11831" />
                    <RANKING order="2" place="2" resultid="12235" />
                    <RANKING order="3" place="3" resultid="12385" />
                    <RANKING order="4" place="4" resultid="12055" />
                    <RANKING order="5" place="5" resultid="11812" />
                    <RANKING order="6" place="6" resultid="12272" />
                    <RANKING order="7" place="7" resultid="12081" />
                    <RANKING order="8" place="8" resultid="12373" />
                    <RANKING order="9" place="9" resultid="12183" />
                    <RANKING order="10" place="10" resultid="11930" />
                    <RANKING order="11" place="11" resultid="12068" />
                    <RANKING order="12" place="12" resultid="11795" />
                    <RANKING order="13" place="-1" resultid="11769" />
                    <RANKING order="14" place="-1" resultid="11893" />
                    <RANKING order="15" place="-1" resultid="12180" />
                    <RANKING order="16" place="-1" resultid="12392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9691" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12020" />
                    <RANKING order="2" place="2" resultid="12032" />
                    <RANKING order="3" place="3" resultid="11840" />
                    <RANKING order="4" place="4" resultid="11818" />
                    <RANKING order="5" place="5" resultid="11837" />
                    <RANKING order="6" place="6" resultid="12222" />
                    <RANKING order="7" place="7" resultid="11823" />
                    <RANKING order="8" place="8" resultid="11950" />
                    <RANKING order="9" place="9" resultid="12104" />
                    <RANKING order="10" place="-1" resultid="12036" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9692" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12048" />
                    <RANKING order="2" place="2" resultid="11999" />
                    <RANKING order="3" place="3" resultid="12573" />
                    <RANKING order="4" place="4" resultid="11808" />
                    <RANKING order="5" place="5" resultid="12363" />
                    <RANKING order="6" place="6" resultid="12170" />
                    <RANKING order="7" place="7" resultid="12398" />
                    <RANKING order="8" place="8" resultid="12132" />
                    <RANKING order="9" place="9" resultid="12633" />
                    <RANKING order="10" place="-1" resultid="11996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9693" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9694" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11880" />
                    <RANKING order="2" place="2" resultid="12023" />
                    <RANKING order="3" place="3" resultid="12502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9695" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12050" />
                    <RANKING order="2" place="2" resultid="12107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9696" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12027" />
                    <RANKING order="2" place="2" resultid="12083" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="9697" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="12961" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12253" />
                    <RANKING order="2" place="2" resultid="11907" />
                    <RANKING order="3" place="3" resultid="11957" />
                    <RANKING order="4" place="4" resultid="12654" />
                    <RANKING order="5" place="5" resultid="12122" />
                    <RANKING order="6" place="6" resultid="12369" />
                    <RANKING order="7" place="7" resultid="12662" />
                    <RANKING order="8" place="8" resultid="12048" />
                    <RANKING order="9" place="9" resultid="11999" />
                    <RANKING order="10" place="9" resultid="12020" />
                    <RANKING order="11" place="11" resultid="12666" />
                    <RANKING order="12" place="12" resultid="12231" />
                    <RANKING order="13" place="13" resultid="11831" />
                    <RANKING order="14" place="14" resultid="12235" />
                    <RANKING order="15" place="15" resultid="12529" />
                    <RANKING order="16" place="16" resultid="12565" />
                    <RANKING order="17" place="17" resultid="12359" />
                    <RANKING order="18" place="18" resultid="12482" />
                    <RANKING order="19" place="19" resultid="12490" />
                    <RANKING order="20" place="20" resultid="12385" />
                    <RANKING order="21" place="21" resultid="12055" />
                    <RANKING order="22" place="22" resultid="12032" />
                    <RANKING order="23" place="23" resultid="11880" />
                    <RANKING order="24" place="24" resultid="12155" />
                    <RANKING order="25" place="25" resultid="11812" />
                    <RANKING order="26" place="26" resultid="12604" />
                    <RANKING order="27" place="27" resultid="12272" />
                    <RANKING order="28" place="28" resultid="12611" />
                    <RANKING order="29" place="29" resultid="12081" />
                    <RANKING order="30" place="30" resultid="11840" />
                    <RANKING order="31" place="31" resultid="12373" />
                    <RANKING order="32" place="32" resultid="12486" />
                    <RANKING order="33" place="33" resultid="12582" />
                    <RANKING order="34" place="34" resultid="11818" />
                    <RANKING order="35" place="35" resultid="12573" />
                    <RANKING order="36" place="36" resultid="12183" />
                    <RANKING order="37" place="37" resultid="11827" />
                    <RANKING order="38" place="38" resultid="12619" />
                    <RANKING order="39" place="39" resultid="11808" />
                    <RANKING order="40" place="40" resultid="11930" />
                    <RANKING order="41" place="41" resultid="12363" />
                    <RANKING order="42" place="42" resultid="12170" />
                    <RANKING order="43" place="43" resultid="12068" />
                    <RANKING order="44" place="44" resultid="12149" />
                    <RANKING order="45" place="45" resultid="11795" />
                    <RANKING order="46" place="46" resultid="11837" />
                    <RANKING order="47" place="47" resultid="12222" />
                    <RANKING order="48" place="48" resultid="11823" />
                    <RANKING order="49" place="49" resultid="12023" />
                    <RANKING order="50" place="50" resultid="12398" />
                    <RANKING order="51" place="51" resultid="12132" />
                    <RANKING order="52" place="52" resultid="12050" />
                    <RANKING order="53" place="53" resultid="11950" />
                    <RANKING order="54" place="54" resultid="12633" />
                    <RANKING order="55" place="55" resultid="12107" />
                    <RANKING order="56" place="56" resultid="12104" />
                    <RANKING order="57" place="57" resultid="12027" />
                    <RANKING order="58" place="58" resultid="12083" />
                    <RANKING order="59" place="59" resultid="12502" />
                    <RANKING order="60" place="-1" resultid="11769" />
                    <RANKING order="61" place="-1" resultid="11996" />
                    <RANKING order="62" place="-1" resultid="12036" />
                    <RANKING order="63" place="-1" resultid="11893" />
                    <RANKING order="64" place="-1" resultid="12180" />
                    <RANKING order="65" place="-1" resultid="12200" />
                    <RANKING order="66" place="-1" resultid="12312" />
                    <RANKING order="67" place="-1" resultid="12377" />
                    <RANKING order="68" place="-1" resultid="12392" />
                    <RANKING order="69" place="-1" resultid="12401" />
                    <RANKING order="70" place="-1" resultid="12420" />
                    <RANKING order="71" place="-1" resultid="12607" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12742" daytime="11:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12743" daytime="11:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12744" daytime="11:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12745" daytime="11:35" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12746" daytime="11:35" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12747" daytime="11:35" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="12748" daytime="11:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="12749" daytime="11:40" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="12805" daytime="11:40" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2164" daytime="11:40" gender="F" number="10" order="10" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10525" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="10526" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="10527" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10528" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12060" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10529" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12177" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10530" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="10531" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12494" />
                    <RANKING order="2" place="2" resultid="12523" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10532" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="10533" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="10534" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="10535" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10536" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10537" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12177" />
                    <RANKING order="2" place="2" resultid="12494" />
                    <RANKING order="3" place="3" resultid="12523" />
                    <RANKING order="4" place="4" resultid="12017" />
                    <RANKING order="5" place="5" resultid="12060" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12750" daytime="11:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2177" daytime="11:45" gender="M" number="11" order="11" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4898" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12140" />
                    <RANKING order="2" place="2" resultid="11791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4899" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12185" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4900" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12670" />
                    <RANKING order="2" place="2" resultid="12525" />
                    <RANKING order="3" place="3" resultid="12285" />
                    <RANKING order="4" place="4" resultid="12440" />
                    <RANKING order="5" place="-1" resultid="12313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4901" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12680" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4902" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12461" />
                    <RANKING order="2" place="2" resultid="12069" />
                    <RANKING order="3" place="-1" resultid="12043" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4903" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12039" />
                    <RANKING order="2" place="2" resultid="12021" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4904" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="4905" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="4906" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="4907" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="4908" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="4909" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="4910" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12140" />
                    <RANKING order="2" place="2" resultid="12039" />
                    <RANKING order="3" place="3" resultid="11791" />
                    <RANKING order="4" place="4" resultid="12670" />
                    <RANKING order="5" place="5" resultid="12525" />
                    <RANKING order="6" place="6" resultid="12285" />
                    <RANKING order="7" place="7" resultid="12680" />
                    <RANKING order="8" place="8" resultid="12021" />
                    <RANKING order="9" place="9" resultid="12185" />
                    <RANKING order="10" place="9" resultid="12461" />
                    <RANKING order="11" place="11" resultid="12440" />
                    <RANKING order="12" place="12" resultid="12069" />
                    <RANKING order="13" place="-1" resultid="12043" />
                    <RANKING order="14" place="-1" resultid="12313" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12751" daytime="11:45" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12752" daytime="11:50" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="10322" daytime="11:50" gender="F" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10323" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="10324" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="10325" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="10326" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="10327" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="10328" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12600" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10329" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10330" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="10331" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="10332" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="10333" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10334" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10335" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12495" />
                    <RANKING order="2" place="2" resultid="12600" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12753" daytime="11:50" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="10336" daytime="11:55" gender="M" number="13" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10337" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10338" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10339" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="10340" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="10341" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="10342" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12224" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10343" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="10344" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10345" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="10346" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="10347" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10348" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10349" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12700" />
                    <RANKING order="2" place="2" resultid="12293" />
                    <RANKING order="3" place="3" resultid="12432" />
                    <RANKING order="4" place="4" resultid="12224" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12754" daytime="11:55" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="10350" daytime="12:00" gender="F" number="14" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10351" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11798" />
                    <RANKING order="2" place="2" resultid="12175" />
                    <RANKING order="3" place="3" resultid="12137" />
                    <RANKING order="4" place="4" resultid="11805" />
                    <RANKING order="5" place="5" resultid="12476" />
                    <RANKING order="6" place="6" resultid="12383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10352" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="10353" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12018" />
                    <RANKING order="2" place="-1" resultid="12507" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10354" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12261" />
                    <RANKING order="2" place="2" resultid="12510" />
                    <RANKING order="3" place="3" resultid="11939" />
                    <RANKING order="4" place="4" resultid="12499" />
                    <RANKING order="5" place="-1" resultid="12218" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10355" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12014" />
                    <RANKING order="2" place="2" resultid="12702" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10356" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12159" />
                    <RANKING order="2" place="2" resultid="12144" />
                    <RANKING order="3" place="3" resultid="12008" />
                    <RANKING order="4" place="4" resultid="12407" />
                    <RANKING order="5" place="5" resultid="12265" />
                    <RANKING order="6" place="6" resultid="12405" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10357" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12247" />
                    <RANKING order="2" place="2" resultid="11896" />
                    <RANKING order="3" place="3" resultid="12243" />
                    <RANKING order="4" place="4" resultid="12298" />
                    <RANKING order="5" place="5" resultid="11802" />
                    <RANKING order="6" place="6" resultid="12098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10358" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11787" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10359" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="10360" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="12011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10361" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10362" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10363" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11798" />
                    <RANKING order="2" place="2" resultid="12261" />
                    <RANKING order="3" place="3" resultid="12175" />
                    <RANKING order="4" place="4" resultid="12247" />
                    <RANKING order="5" place="5" resultid="12159" />
                    <RANKING order="6" place="6" resultid="12014" />
                    <RANKING order="7" place="7" resultid="12510" />
                    <RANKING order="8" place="8" resultid="11896" />
                    <RANKING order="9" place="9" resultid="12243" />
                    <RANKING order="10" place="10" resultid="12137" />
                    <RANKING order="11" place="11" resultid="12298" />
                    <RANKING order="12" place="12" resultid="11805" />
                    <RANKING order="13" place="13" resultid="12144" />
                    <RANKING order="14" place="14" resultid="12008" />
                    <RANKING order="15" place="15" resultid="12702" />
                    <RANKING order="16" place="16" resultid="11802" />
                    <RANKING order="17" place="17" resultid="12018" />
                    <RANKING order="18" place="17" resultid="12407" />
                    <RANKING order="19" place="19" resultid="12098" />
                    <RANKING order="20" place="20" resultid="11939" />
                    <RANKING order="21" place="21" resultid="12265" />
                    <RANKING order="22" place="22" resultid="12476" />
                    <RANKING order="23" place="23" resultid="12499" />
                    <RANKING order="24" place="24" resultid="11787" />
                    <RANKING order="25" place="25" resultid="12383" />
                    <RANKING order="26" place="26" resultid="12405" />
                    <RANKING order="27" place="-1" resultid="12507" />
                    <RANKING order="28" place="-1" resultid="12011" />
                    <RANKING order="29" place="-1" resultid="12218" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12755" daytime="12:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12756" daytime="12:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12757" daytime="12:05" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12806" daytime="12:05" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="10364" daytime="12:05" gender="M" number="15" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10365" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11792" />
                    <RANKING order="2" place="2" resultid="11778" />
                    <RANKING order="3" place="3" resultid="12352" />
                    <RANKING order="4" place="4" resultid="12228" />
                    <RANKING order="5" place="5" resultid="12232" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10366" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12667" />
                    <RANKING order="2" place="2" resultid="11915" />
                    <RANKING order="3" place="3" resultid="12491" />
                    <RANKING order="4" place="-1" resultid="12421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10367" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12526" />
                    <RANKING order="2" place="2" resultid="12650" />
                    <RANKING order="3" place="3" resultid="12664" />
                    <RANKING order="4" place="4" resultid="12156" />
                    <RANKING order="5" place="5" resultid="12441" />
                    <RANKING order="6" place="6" resultid="12147" />
                    <RANKING order="7" place="-1" resultid="12426" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10368" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12459" />
                    <RANKING order="2" place="2" resultid="12530" />
                    <RANKING order="3" place="3" resultid="12566" />
                    <RANKING order="4" place="4" resultid="12605" />
                    <RANKING order="5" place="5" resultid="12620" />
                    <RANKING order="6" place="6" resultid="11828" />
                    <RANKING order="7" place="-1" resultid="12378" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10369" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12636" />
                    <RANKING order="2" place="2" resultid="12273" />
                    <RANKING order="3" place="3" resultid="12071" />
                    <RANKING order="4" place="4" resultid="12386" />
                    <RANKING order="5" place="5" resultid="11832" />
                    <RANKING order="6" place="6" resultid="11931" />
                    <RANKING order="7" place="-1" resultid="11770" />
                    <RANKING order="8" place="-1" resultid="12181" />
                    <RANKING order="9" place="-1" resultid="12393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10370" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12319" />
                    <RANKING order="2" place="2" resultid="11841" />
                    <RANKING order="3" place="3" resultid="11834" />
                    <RANKING order="4" place="4" resultid="11824" />
                    <RANKING order="5" place="5" resultid="11838" />
                    <RANKING order="6" place="6" resultid="12105" />
                    <RANKING order="7" place="7" resultid="11951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10371" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12000" />
                    <RANKING order="2" place="2" resultid="12171" />
                    <RANKING order="3" place="3" resultid="11809" />
                    <RANKING order="4" place="4" resultid="12640" />
                    <RANKING order="5" place="5" resultid="12574" />
                    <RANKING order="6" place="6" resultid="12364" />
                    <RANKING order="7" place="7" resultid="12323" />
                    <RANKING order="8" place="8" resultid="12133" />
                    <RANKING order="9" place="9" resultid="12634" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10372" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12003" />
                    <RANKING order="2" place="2" resultid="12250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10373" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12472" />
                    <RANKING order="2" place="2" resultid="12024" />
                    <RANKING order="3" place="3" resultid="12075" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10374" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12051" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10375" agemax="79" agemin="75">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12084" />
                    <RANKING order="2" place="2" resultid="12028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10376" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10377" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11792" />
                    <RANKING order="2" place="1" resultid="12003" />
                    <RANKING order="3" place="3" resultid="12526" />
                    <RANKING order="4" place="4" resultid="11778" />
                    <RANKING order="5" place="5" resultid="12000" />
                    <RANKING order="6" place="6" resultid="12650" />
                    <RANKING order="7" place="7" resultid="12664" />
                    <RANKING order="8" place="8" resultid="12352" />
                    <RANKING order="9" place="9" resultid="12636" />
                    <RANKING order="10" place="10" resultid="12319" />
                    <RANKING order="11" place="11" resultid="12459" />
                    <RANKING order="12" place="12" resultid="12472" />
                    <RANKING order="13" place="13" resultid="12667" />
                    <RANKING order="14" place="14" resultid="12228" />
                    <RANKING order="15" place="15" resultid="12530" />
                    <RANKING order="16" place="16" resultid="12024" />
                    <RANKING order="17" place="17" resultid="12566" />
                    <RANKING order="18" place="18" resultid="11915" />
                    <RANKING order="19" place="19" resultid="12273" />
                    <RANKING order="20" place="20" resultid="11841" />
                    <RANKING order="21" place="21" resultid="11834" />
                    <RANKING order="22" place="22" resultid="12071" />
                    <RANKING order="23" place="23" resultid="12171" />
                    <RANKING order="24" place="24" resultid="11809" />
                    <RANKING order="25" place="25" resultid="12232" />
                    <RANKING order="26" place="26" resultid="12605" />
                    <RANKING order="27" place="27" resultid="12386" />
                    <RANKING order="28" place="28" resultid="12640" />
                    <RANKING order="29" place="29" resultid="12574" />
                    <RANKING order="30" place="30" resultid="11832" />
                    <RANKING order="31" place="31" resultid="12084" />
                    <RANKING order="32" place="32" resultid="12364" />
                    <RANKING order="33" place="33" resultid="12620" />
                    <RANKING order="34" place="34" resultid="11824" />
                    <RANKING order="35" place="35" resultid="11838" />
                    <RANKING order="36" place="36" resultid="11828" />
                    <RANKING order="37" place="37" resultid="12051" />
                    <RANKING order="38" place="38" resultid="12156" />
                    <RANKING order="39" place="39" resultid="12491" />
                    <RANKING order="40" place="40" resultid="11931" />
                    <RANKING order="41" place="41" resultid="12250" />
                    <RANKING order="42" place="42" resultid="12323" />
                    <RANKING order="43" place="43" resultid="12028" />
                    <RANKING order="44" place="44" resultid="12133" />
                    <RANKING order="45" place="45" resultid="12441" />
                    <RANKING order="46" place="46" resultid="12105" />
                    <RANKING order="47" place="47" resultid="12075" />
                    <RANKING order="48" place="48" resultid="12147" />
                    <RANKING order="49" place="49" resultid="12634" />
                    <RANKING order="50" place="50" resultid="11951" />
                    <RANKING order="51" place="-1" resultid="12426" />
                    <RANKING order="52" place="-1" resultid="11770" />
                    <RANKING order="53" place="-1" resultid="12181" />
                    <RANKING order="54" place="-1" resultid="12378" />
                    <RANKING order="55" place="-1" resultid="12393" />
                    <RANKING order="56" place="-1" resultid="12421" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12758" daytime="12:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12759" daytime="12:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12760" daytime="12:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12761" daytime="12:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12762" daytime="12:15" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12763" daytime="12:15" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="12807" daytime="12:15" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1061" daytime="12:30" gender="X" number="16" order="17" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="EUR" value="350" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2103" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11845" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2104" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12334" />
                    <RANKING order="2" place="2" resultid="12208" />
                    <RANKING order="3" place="-1" resultid="12412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2105" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12532" />
                    <RANKING order="2" place="2" resultid="12338" />
                    <RANKING order="3" place="3" resultid="12090" />
                    <RANKING order="4" place="4" resultid="12643" />
                    <RANKING order="5" place="5" resultid="12413" />
                    <RANKING order="6" place="-1" resultid="12207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2106" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12342" />
                    <RANKING order="2" place="-1" resultid="12093" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2107" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="2108" agemax="319" agemin="280" calculate="TOTAL" />
                <AGEGROUP agegroupid="2109" agemax="359" agemin="320" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12764" daytime="12:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12765" daytime="12:35" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2021-12-04" daytime="15:00" endtime="17:31" name="2ª Jornada" number="2" warmupfrom="14:00" warmupuntil="14:45">
          <EVENTS>
            <EVENT eventid="10378" daytime="15:00" gender="X" number="17" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="EUR" value="350" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10379" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10380" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11990" />
                    <RANKING order="2" place="2" resultid="12339" />
                    <RANKING order="3" place="3" resultid="12531" />
                    <RANKING order="4" place="4" resultid="12454" />
                    <RANKING order="5" place="-1" resultid="12205" />
                    <RANKING order="6" place="-1" resultid="12411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10381" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12341" />
                    <RANKING order="2" place="2" resultid="12644" />
                    <RANKING order="3" place="3" resultid="12692" />
                    <RANKING order="4" place="4" resultid="11844" />
                    <RANKING order="5" place="5" resultid="12942" />
                    <RANKING order="6" place="6" resultid="11953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10382" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12583" />
                    <RANKING order="2" place="2" resultid="12558" />
                    <RANKING order="3" place="3" resultid="12346" />
                    <RANKING order="4" place="4" resultid="12416" />
                    <RANKING order="5" place="5" resultid="12206" />
                    <RANKING order="6" place="6" resultid="11843" />
                    <RANKING order="7" place="-1" resultid="12091" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10383" agemax="279" agemin="240" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12535" />
                    <RANKING order="2" place="2" resultid="12349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10384" agemax="319" agemin="280" calculate="TOTAL" />
                <AGEGROUP agegroupid="10385" agemax="359" agemin="320" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12766" daytime="15:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12767" daytime="15:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12768" daytime="15:10" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1118" daytime="15:10" gender="F" number="18" order="2" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4846" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4847" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12327" />
                    <RANKING order="2" place="2" resultid="12192" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4848" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="4849" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12166" />
                    <RANKING order="2" place="2" resultid="12130" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4850" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="4851" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="4852" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="4853" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="4854" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="4855" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="4856" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="4857" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="4858" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11761" />
                    <RANKING order="2" place="2" resultid="12166" />
                    <RANKING order="3" place="3" resultid="12130" />
                    <RANKING order="4" place="4" resultid="12327" />
                    <RANKING order="5" place="5" resultid="12192" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12769" daytime="15:10" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="10455">
                  <FEE currency="EUR" value="400" />
                </TIMESTANDARDREF>
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1131" daytime="15:20" gender="M" number="19" order="3" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4924" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="4925" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4926" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12118" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4927" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="4928" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4929" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12480" />
                    <RANKING order="2" place="2" resultid="12040" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4930" agemax="59" agemin="55" />
                <AGEGROUP agegroupid="4931" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="4932" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="4933" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="4934" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="4935" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="4936" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12480" />
                    <RANKING order="2" place="2" resultid="12040" />
                    <RANKING order="3" place="3" resultid="12517" />
                    <RANKING order="4" place="4" resultid="12118" />
                    <RANKING order="5" place="5" resultid="12433" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12770" daytime="15:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="10441">
                  <FEE currency="EUR" value="400" />
                </TIMESTANDARDREF>
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="9711" daytime="15:25" gender="F" number="20" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10551" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12659" />
                    <RANKING order="2" place="2" resultid="12423" />
                    <RANKING order="3" place="3" resultid="12428" />
                    <RANKING order="4" place="4" resultid="12382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10552" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12316" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10553" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12258" />
                    <RANKING order="2" place="2" resultid="12152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10554" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12677" />
                    <RANKING order="2" place="2" resultid="12269" />
                    <RANKING order="3" place="3" resultid="12579" />
                    <RANKING order="4" place="4" resultid="11856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10555" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12703" />
                    <RANKING order="2" place="-1" resultid="11993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10556" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12601" />
                    <RANKING order="2" place="2" resultid="12160" />
                    <RANKING order="3" place="3" resultid="12550" />
                    <RANKING order="4" place="4" resultid="12408" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10557" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10558" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10559" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="10560" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="10561" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10562" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10563" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12659" />
                    <RANKING order="2" place="2" resultid="12677" />
                    <RANKING order="3" place="3" resultid="12258" />
                    <RANKING order="4" place="4" resultid="12269" />
                    <RANKING order="5" place="5" resultid="12423" />
                    <RANKING order="6" place="6" resultid="12579" />
                    <RANKING order="7" place="7" resultid="12428" />
                    <RANKING order="8" place="8" resultid="12152" />
                    <RANKING order="9" place="9" resultid="12601" />
                    <RANKING order="10" place="10" resultid="12160" />
                    <RANKING order="11" place="11" resultid="12703" />
                    <RANKING order="12" place="12" resultid="12276" />
                    <RANKING order="13" place="13" resultid="12550" />
                    <RANKING order="14" place="14" resultid="12408" />
                    <RANKING order="15" place="15" resultid="12316" />
                    <RANKING order="16" place="16" resultid="12382" />
                    <RANKING order="17" place="17" resultid="11856" />
                    <RANKING order="18" place="18" resultid="12198" />
                    <RANKING order="19" place="-1" resultid="11993" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12771" daytime="15:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12772" daytime="15:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12808" daytime="15:35" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="9737" daytime="15:35" gender="M" number="21" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10590" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11779" />
                    <RANKING order="2" place="2" resultid="12294" />
                    <RANKING order="3" place="3" resultid="12655" />
                    <RANKING order="4" place="4" resultid="12370" />
                    <RANKING order="5" place="5" resultid="11947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10591" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12254" />
                    <RANKING order="2" place="2" resultid="11908" />
                    <RANKING order="3" place="3" resultid="12668" />
                    <RANKING order="4" place="4" resultid="12492" />
                    <RANKING order="5" place="5" resultid="12451" />
                    <RANKING order="6" place="-1" resultid="12201" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10592" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12663" />
                    <RANKING order="2" place="2" resultid="11875" />
                    <RANKING order="3" place="3" resultid="12064" />
                    <RANKING order="4" place="4" resultid="12148" />
                    <RANKING order="5" place="-1" resultid="12608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10593" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11958" />
                    <RANKING order="2" place="2" resultid="11867" />
                    <RANKING order="3" place="3" resultid="12612" />
                    <RANKING order="4" place="4" resultid="12621" />
                    <RANKING order="5" place="5" resultid="12447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10594" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12468" />
                    <RANKING order="2" place="2" resultid="12236" />
                    <RANKING order="3" place="3" resultid="12462" />
                    <RANKING order="4" place="4" resultid="11862" />
                    <RANKING order="5" place="5" resultid="12374" />
                    <RANKING order="6" place="6" resultid="11796" />
                    <RANKING order="7" place="7" resultid="11943" />
                    <RANKING order="8" place="8" resultid="12437" />
                    <RANKING order="9" place="-1" resultid="11774" />
                    <RANKING order="10" place="-1" resultid="12110" />
                    <RANKING order="11" place="-1" resultid="12615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10595" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11842" />
                    <RANKING order="2" place="2" resultid="11869" />
                    <RANKING order="3" place="3" resultid="12444" />
                    <RANKING order="4" place="4" resultid="12126" />
                    <RANKING order="5" place="5" resultid="12539" />
                    <RANKING order="6" place="6" resultid="11952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10596" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12290" />
                    <RANKING order="2" place="2" resultid="12543" />
                    <RANKING order="3" place="3" resultid="12365" />
                    <RANKING order="4" place="4" resultid="12399" />
                    <RANKING order="5" place="5" resultid="12635" />
                    <RANKING order="6" place="-1" resultid="11872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10597" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="10598" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12569" />
                    <RANKING order="2" place="2" resultid="12076" />
                    <RANKING order="3" place="3" resultid="12503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10599" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10600" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10601" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10602" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11958" />
                    <RANKING order="2" place="2" resultid="11779" />
                    <RANKING order="3" place="3" resultid="12254" />
                    <RANKING order="4" place="4" resultid="12294" />
                    <RANKING order="5" place="5" resultid="12663" />
                    <RANKING order="6" place="6" resultid="11908" />
                    <RANKING order="7" place="7" resultid="12655" />
                    <RANKING order="8" place="8" resultid="12370" />
                    <RANKING order="9" place="9" resultid="12468" />
                    <RANKING order="10" place="9" resultid="12290" />
                    <RANKING order="11" place="11" resultid="12236" />
                    <RANKING order="12" place="12" resultid="11867" />
                    <RANKING order="13" place="13" resultid="12668" />
                    <RANKING order="14" place="14" resultid="12462" />
                    <RANKING order="15" place="15" resultid="12569" />
                    <RANKING order="16" place="16" resultid="12543" />
                    <RANKING order="17" place="17" resultid="11875" />
                    <RANKING order="18" place="18" resultid="11862" />
                    <RANKING order="19" place="19" resultid="12365" />
                    <RANKING order="20" place="20" resultid="12492" />
                    <RANKING order="21" place="21" resultid="11842" />
                    <RANKING order="22" place="22" resultid="11869" />
                    <RANKING order="23" place="23" resultid="12451" />
                    <RANKING order="24" place="23" resultid="12612" />
                    <RANKING order="25" place="25" resultid="12374" />
                    <RANKING order="26" place="26" resultid="11947" />
                    <RANKING order="27" place="27" resultid="12561" />
                    <RANKING order="28" place="28" resultid="12444" />
                    <RANKING order="29" place="29" resultid="12126" />
                    <RANKING order="30" place="30" resultid="12539" />
                    <RANKING order="31" place="31" resultid="12064" />
                    <RANKING order="32" place="32" resultid="11796" />
                    <RANKING order="33" place="33" resultid="12148" />
                    <RANKING order="34" place="34" resultid="11943" />
                    <RANKING order="35" place="35" resultid="12621" />
                    <RANKING order="36" place="36" resultid="12437" />
                    <RANKING order="37" place="37" resultid="12399" />
                    <RANKING order="38" place="38" resultid="12076" />
                    <RANKING order="39" place="39" resultid="12447" />
                    <RANKING order="40" place="40" resultid="12635" />
                    <RANKING order="41" place="41" resultid="11952" />
                    <RANKING order="42" place="42" resultid="12503" />
                    <RANKING order="43" place="-1" resultid="11774" />
                    <RANKING order="44" place="-1" resultid="12110" />
                    <RANKING order="45" place="-1" resultid="11872" />
                    <RANKING order="46" place="-1" resultid="12201" />
                    <RANKING order="47" place="-1" resultid="12608" />
                    <RANKING order="48" place="-1" resultid="12615" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12773" daytime="15:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12774" daytime="15:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12775" daytime="15:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12776" daytime="15:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12777" daytime="15:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="12809" daytime="15:50" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1144" daytime="15:50" gender="F" number="22" order="6" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4859" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12632" />
                    <RANKING order="2" place="2" resultid="12685" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4860" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="4861" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12259" />
                    <RANKING order="2" place="2" resultid="12153" />
                    <RANKING order="3" place="3" resultid="11935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4862" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12630" />
                    <RANKING order="2" place="2" resultid="12547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4863" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="4864" agemax="54" agemin="50" />
                <AGEGROUP agegroupid="4865" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12239" />
                    <RANKING order="2" place="2" resultid="12244" />
                    <RANKING order="3" place="3" resultid="12299" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4866" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="4867" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="4868" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="4869" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="4870" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="4871" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12632" />
                    <RANKING order="2" place="2" resultid="12259" />
                    <RANKING order="3" place="3" resultid="12239" />
                    <RANKING order="4" place="4" resultid="12244" />
                    <RANKING order="5" place="5" resultid="12153" />
                    <RANKING order="6" place="6" resultid="12299" />
                    <RANKING order="7" place="7" resultid="12630" />
                    <RANKING order="8" place="8" resultid="12547" />
                    <RANKING order="9" place="9" resultid="11935" />
                    <RANKING order="10" place="10" resultid="12685" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12778" daytime="15:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12810" daytime="15:55" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1157" daytime="16:00" gender="M" number="23" order="7" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5521" agemax="29" agemin="25" />
                <AGEGROUP agegroupid="5522" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12112" />
                    <RANKING order="2" place="2" resultid="12123" />
                    <RANKING order="3" place="3" resultid="12186" />
                    <RANKING order="4" place="4" resultid="11916" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5523" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12672" />
                    <RANKING order="2" place="2" resultid="12286" />
                    <RANKING order="3" place="3" resultid="12442" />
                    <RANKING order="4" place="4" resultid="12487" />
                    <RANKING order="5" place="5" resultid="12065" />
                    <RANKING order="6" place="6" resultid="12355" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5524" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11959" />
                    <RANKING order="2" place="2" resultid="12567" />
                    <RANKING order="3" place="3" resultid="12115" />
                    <RANKING order="4" place="4" resultid="12357" />
                    <RANKING order="5" place="-1" resultid="12681" />
                    <RANKING order="6" place="-1" resultid="12379" />
                    <RANKING order="7" place="-1" resultid="12402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5525" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12518" />
                    <RANKING order="2" place="2" resultid="12282" />
                    <RANKING order="3" place="3" resultid="12304" />
                    <RANKING order="4" place="4" resultid="12469" />
                    <RANKING order="5" place="5" resultid="11863" />
                    <RANKING order="6" place="6" resultid="12101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5526" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12367" />
                    <RANKING order="2" place="2" resultid="11859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5527" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12553" />
                    <RANKING order="2" place="2" resultid="12302" />
                    <RANKING order="3" place="3" resultid="11997" />
                    <RANKING order="4" place="4" resultid="12575" />
                    <RANKING order="5" place="5" resultid="12639" />
                    <RANKING order="6" place="6" resultid="12515" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5528" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11888" />
                    <RANKING order="2" place="2" resultid="12483" />
                    <RANKING order="3" place="3" resultid="12251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5529" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11881" />
                    <RANKING order="2" place="2" resultid="12570" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5530" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="5531" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="5532" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="5533" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11888" />
                    <RANKING order="2" place="2" resultid="11881" />
                    <RANKING order="3" place="3" resultid="12672" />
                    <RANKING order="4" place="4" resultid="12518" />
                    <RANKING order="5" place="5" resultid="11959" />
                    <RANKING order="6" place="6" resultid="12286" />
                    <RANKING order="7" place="7" resultid="12112" />
                    <RANKING order="8" place="8" resultid="12123" />
                    <RANKING order="9" place="9" resultid="12553" />
                    <RANKING order="10" place="10" resultid="12302" />
                    <RANKING order="11" place="11" resultid="12483" />
                    <RANKING order="12" place="12" resultid="12282" />
                    <RANKING order="13" place="13" resultid="12567" />
                    <RANKING order="14" place="14" resultid="12304" />
                    <RANKING order="15" place="15" resultid="12186" />
                    <RANKING order="16" place="16" resultid="12570" />
                    <RANKING order="17" place="17" resultid="12469" />
                    <RANKING order="18" place="18" resultid="12367" />
                    <RANKING order="19" place="19" resultid="12115" />
                    <RANKING order="20" place="20" resultid="11997" />
                    <RANKING order="21" place="21" resultid="11859" />
                    <RANKING order="22" place="22" resultid="11916" />
                    <RANKING order="23" place="23" resultid="12251" />
                    <RANKING order="24" place="24" resultid="12575" />
                    <RANKING order="25" place="25" resultid="11863" />
                    <RANKING order="26" place="26" resultid="12442" />
                    <RANKING order="27" place="27" resultid="12101" />
                    <RANKING order="28" place="28" resultid="12487" />
                    <RANKING order="29" place="29" resultid="12639" />
                    <RANKING order="30" place="30" resultid="12357" />
                    <RANKING order="31" place="31" resultid="12515" />
                    <RANKING order="32" place="32" resultid="12065" />
                    <RANKING order="33" place="33" resultid="12355" />
                    <RANKING order="34" place="-1" resultid="12681" />
                    <RANKING order="35" place="-1" resultid="12379" />
                    <RANKING order="36" place="-1" resultid="12402" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12779" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12780" daytime="16:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12781" daytime="16:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12782" daytime="16:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12811" daytime="16:20" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="10386" daytime="16:20" gender="F" number="24" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10564" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12648" />
                    <RANKING order="2" place="2" resultid="12477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10565" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12329" />
                    <RANKING order="2" place="2" resultid="12317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10566" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12332" />
                    <RANKING order="2" place="2" resultid="12508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10567" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12500" />
                    <RANKING order="2" place="2" resultid="12629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10568" agemax="49" agemin="45" />
                <AGEGROUP agegroupid="10569" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12465" />
                    <RANKING order="2" place="2" resultid="12551" />
                    <RANKING order="3" place="3" resultid="12690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10570" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11852" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10571" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12309" />
                    <RANKING order="2" place="2" resultid="12277" />
                    <RANKING order="3" place="3" resultid="12195" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10572" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="10573" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="10574" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10575" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10576" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12329" />
                    <RANKING order="2" place="2" resultid="11852" />
                    <RANKING order="3" place="3" resultid="12648" />
                    <RANKING order="4" place="4" resultid="12465" />
                    <RANKING order="5" place="5" resultid="12332" />
                    <RANKING order="6" place="6" resultid="12477" />
                    <RANKING order="7" place="7" resultid="12309" />
                    <RANKING order="8" place="8" resultid="12500" />
                    <RANKING order="9" place="9" resultid="12629" />
                    <RANKING order="10" place="10" resultid="12551" />
                    <RANKING order="11" place="11" resultid="12317" />
                    <RANKING order="12" place="11" resultid="12277" />
                    <RANKING order="13" place="13" resultid="12195" />
                    <RANKING order="14" place="14" resultid="12508" />
                    <RANKING order="15" place="15" resultid="12690" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12783" daytime="16:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12784" daytime="16:25" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="10399" daytime="16:30" gender="M" number="25" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10603" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10604" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="10605" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10606" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="10607" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="11771" />
                    <RANKING order="2" place="-1" resultid="12556" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10608" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10609" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12554" />
                    <RANKING order="2" place="2" resultid="12544" />
                    <RANKING order="3" place="3" resultid="12324" />
                    <RANKING order="4" place="-1" resultid="12688" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10610" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="10611" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12025" />
                    <RANKING order="2" place="-1" resultid="12473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10612" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="10613" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10614" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10615" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12360" />
                    <RANKING order="2" place="2" resultid="12025" />
                    <RANKING order="3" place="3" resultid="12554" />
                    <RANKING order="4" place="4" resultid="11874" />
                    <RANKING order="5" place="5" resultid="12544" />
                    <RANKING order="6" place="6" resultid="12540" />
                    <RANKING order="7" place="7" resultid="12324" />
                    <RANKING order="8" place="-1" resultid="12473" />
                    <RANKING order="9" place="-1" resultid="12688" />
                    <RANKING order="10" place="-1" resultid="11771" />
                    <RANKING order="11" place="-1" resultid="12556" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12785" daytime="16:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12786" daytime="16:30" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="9763" daytime="16:35" gender="F" number="26" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10577" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11799" />
                    <RANKING order="2" place="2" resultid="11806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10578" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="10579" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12331" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10580" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12678" />
                    <RANKING order="2" place="2" resultid="11821" />
                    <RANKING order="3" place="3" resultid="12548" />
                    <RANKING order="4" place="4" resultid="11940" />
                    <RANKING order="5" place="5" resultid="11857" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10581" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12178" />
                    <RANKING order="2" place="-1" resultid="11994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10582" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12145" />
                    <RANKING order="2" place="2" resultid="12409" />
                    <RANKING order="3" place="3" resultid="12266" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10583" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12240" />
                    <RANKING order="2" place="2" resultid="12245" />
                    <RANKING order="3" place="3" resultid="11803" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10584" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="10585" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="10586" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="10587" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10588" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10589" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11799" />
                    <RANKING order="2" place="2" resultid="12240" />
                    <RANKING order="3" place="3" resultid="12678" />
                    <RANKING order="4" place="4" resultid="12245" />
                    <RANKING order="5" place="5" resultid="12178" />
                    <RANKING order="6" place="6" resultid="11806" />
                    <RANKING order="7" place="7" resultid="11821" />
                    <RANKING order="8" place="8" resultid="12145" />
                    <RANKING order="9" place="9" resultid="12409" />
                    <RANKING order="10" place="10" resultid="12548" />
                    <RANKING order="11" place="11" resultid="12331" />
                    <RANKING order="12" place="11" resultid="12266" />
                    <RANKING order="13" place="13" resultid="11940" />
                    <RANKING order="14" place="14" resultid="11803" />
                    <RANKING order="15" place="15" resultid="11857" />
                    <RANKING order="16" place="-1" resultid="11994" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12787" daytime="16:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12788" daytime="16:35" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="9789" daytime="16:40" gender="M" number="27" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10616" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12353" />
                    <RANKING order="2" place="2" resultid="11793" />
                    <RANKING order="3" place="3" resultid="11948" />
                    <RANKING order="4" place="4" resultid="12233" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10617" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12699" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10618" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12527" />
                    <RANKING order="2" place="2" resultid="12651" />
                    <RANKING order="3" place="3" resultid="12488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10619" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11866" />
                    <RANKING order="2" place="2" resultid="12613" />
                    <RANKING order="3" place="3" resultid="11829" />
                    <RANKING order="4" place="4" resultid="12448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10620" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11813" />
                    <RANKING order="2" place="2" resultid="12390" />
                    <RANKING order="3" place="3" resultid="12438" />
                    <RANKING order="4" place="4" resultid="11944" />
                    <RANKING order="5" place="-1" resultid="12557" />
                    <RANKING order="6" place="-1" resultid="12616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10621" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12320" />
                    <RANKING order="2" place="2" resultid="11860" />
                    <RANKING order="3" place="3" resultid="12225" />
                    <RANKING order="4" place="4" resultid="11825" />
                    <RANKING order="5" place="5" resultid="12445" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10622" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12001" />
                    <RANKING order="2" place="2" resultid="12172" />
                    <RANKING order="3" place="3" resultid="11810" />
                    <RANKING order="4" place="4" resultid="12325" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10623" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12004" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10624" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="10625" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10626" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10627" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10628" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12004" />
                    <RANKING order="2" place="2" resultid="12353" />
                    <RANKING order="3" place="3" resultid="12001" />
                    <RANKING order="4" place="4" resultid="12527" />
                    <RANKING order="5" place="5" resultid="11793" />
                    <RANKING order="6" place="6" resultid="12651" />
                    <RANKING order="7" place="7" resultid="12699" />
                    <RANKING order="8" place="8" resultid="12320" />
                    <RANKING order="9" place="9" resultid="11860" />
                    <RANKING order="10" place="10" resultid="11866" />
                    <RANKING order="11" place="10" resultid="12172" />
                    <RANKING order="12" place="12" resultid="12562" />
                    <RANKING order="13" place="13" resultid="11813" />
                    <RANKING order="14" place="14" resultid="12613" />
                    <RANKING order="15" place="15" resultid="11810" />
                    <RANKING order="16" place="16" resultid="11948" />
                    <RANKING order="17" place="17" resultid="12225" />
                    <RANKING order="18" place="18" resultid="12233" />
                    <RANKING order="19" place="19" resultid="12390" />
                    <RANKING order="20" place="20" resultid="11825" />
                    <RANKING order="21" place="21" resultid="12445" />
                    <RANKING order="22" place="22" resultid="11829" />
                    <RANKING order="23" place="23" resultid="12488" />
                    <RANKING order="24" place="24" resultid="12325" />
                    <RANKING order="25" place="25" resultid="12448" />
                    <RANKING order="26" place="26" resultid="12438" />
                    <RANKING order="27" place="27" resultid="11944" />
                    <RANKING order="28" place="-1" resultid="12557" />
                    <RANKING order="29" place="-1" resultid="12616" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12789" daytime="16:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12790" daytime="16:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12791" daytime="16:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12812" daytime="16:45" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2190" daytime="16:50" gender="F" number="28" order="12" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4872" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11762" />
                    <RANKING order="2" place="2" resultid="12424" />
                    <RANKING order="3" place="3" resultid="12429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4873" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="4874" agemax="39" agemin="35" />
                <AGEGROUP agegroupid="4875" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12167" />
                    <RANKING order="2" place="2" resultid="12511" />
                    <RANKING order="3" place="3" resultid="12580" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4876" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12015" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4877" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12161" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4878" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4879" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12278" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4880" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="4881" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="4882" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="4883" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="4884" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11762" />
                    <RANKING order="2" place="2" resultid="12167" />
                    <RANKING order="3" place="3" resultid="12424" />
                    <RANKING order="4" place="4" resultid="12511" />
                    <RANKING order="5" place="5" resultid="12015" />
                    <RANKING order="6" place="6" resultid="12161" />
                    <RANKING order="7" place="7" resultid="12429" />
                    <RANKING order="8" place="8" resultid="12580" />
                    <RANKING order="9" place="9" resultid="12099" />
                    <RANKING order="10" place="10" resultid="12278" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12792" daytime="16:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12813" daytime="16:55" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2203" daytime="17:00" gender="M" number="29" order="13" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4911" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12141" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4912" agemax="34" agemin="30" />
                <AGEGROUP agegroupid="4913" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12652" />
                    <RANKING order="2" place="2" resultid="11876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4914" agemax="44" agemin="40" />
                <AGEGROUP agegroupid="4915" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12305" />
                    <RANKING order="2" place="2" resultid="11932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4916" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12321" />
                    <RANKING order="2" place="2" resultid="11835" />
                    <RANKING order="3" place="3" resultid="12226" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4917" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12545" />
                    <RANKING order="2" place="2" resultid="12134" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4918" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="4919" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12571" />
                    <RANKING order="2" place="-1" resultid="12504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4920" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12108" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4921" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="4922" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="4923" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12141" />
                    <RANKING order="2" place="2" resultid="12652" />
                    <RANKING order="3" place="3" resultid="12305" />
                    <RANKING order="4" place="4" resultid="12321" />
                    <RANKING order="5" place="5" resultid="11835" />
                    <RANKING order="6" place="6" resultid="11876" />
                    <RANKING order="7" place="7" resultid="12545" />
                    <RANKING order="8" place="8" resultid="12226" />
                    <RANKING order="9" place="9" resultid="11932" />
                    <RANKING order="10" place="10" resultid="12571" />
                    <RANKING order="11" place="11" resultid="12108" />
                    <RANKING order="12" place="12" resultid="12134" />
                    <RANKING order="13" place="-1" resultid="12504" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12793" daytime="17:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12794" daytime="17:05" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="10412" daytime="17:10" gender="F" number="30" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10413" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12660" />
                    <RANKING order="2" place="2" resultid="12686" />
                    <RANKING order="3" place="-1" resultid="11763" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10414" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12328" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10415" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11936" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10416" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12262" />
                    <RANKING order="2" place="2" resultid="12512" />
                    <RANKING order="3" place="3" resultid="12270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10417" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12216" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10418" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10419" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11853" />
                    <RANKING order="2" place="2" resultid="12496" />
                    <RANKING order="3" place="3" resultid="12241" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10420" agemax="64" agemin="60" />
                <AGEGROUP agegroupid="10421" agemax="69" agemin="65" />
                <AGEGROUP agegroupid="10422" agemax="74" agemin="70" />
                <AGEGROUP agegroupid="10423" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10424" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10425" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12328" />
                    <RANKING order="2" place="2" resultid="12660" />
                    <RANKING order="3" place="3" resultid="12262" />
                    <RANKING order="4" place="4" resultid="12216" />
                    <RANKING order="5" place="5" resultid="12512" />
                    <RANKING order="6" place="6" resultid="12270" />
                    <RANKING order="7" place="7" resultid="11853" />
                    <RANKING order="8" place="8" resultid="12496" />
                    <RANKING order="9" place="9" resultid="11936" />
                    <RANKING order="10" place="10" resultid="12241" />
                    <RANKING order="11" place="11" resultid="12602" />
                    <RANKING order="12" place="12" resultid="12686" />
                    <RANKING order="13" place="-1" resultid="11763" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12795" daytime="17:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12796" daytime="17:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="10426" daytime="17:15" gender="M" number="31" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="EUR" value="300" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="10427" agemax="29" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12295" />
                    <RANKING order="2" place="2" resultid="11780" />
                    <RANKING order="3" place="3" resultid="12656" />
                    <RANKING order="4" place="4" resultid="12361" />
                    <RANKING order="5" place="5" resultid="12229" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10428" agemax="34" agemin="30">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12255" />
                    <RANKING order="2" place="2" resultid="11909" />
                    <RANKING order="3" place="3" resultid="12124" />
                    <RANKING order="4" place="4" resultid="12113" />
                    <RANKING order="5" place="-1" resultid="12452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10429" agemax="39" agemin="35">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12287" />
                    <RANKING order="2" place="2" resultid="12157" />
                    <RANKING order="3" place="3" resultid="12066" />
                    <RANKING order="4" place="-1" resultid="12609" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10430" agemax="44" agemin="40">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12682" />
                    <RANKING order="2" place="2" resultid="12116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10431" agemax="49" agemin="45">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12519" />
                    <RANKING order="2" place="2" resultid="12637" />
                    <RANKING order="3" place="3" resultid="12306" />
                    <RANKING order="4" place="4" resultid="12237" />
                    <RANKING order="5" place="5" resultid="12463" />
                    <RANKING order="6" place="6" resultid="11814" />
                    <RANKING order="7" place="7" resultid="12283" />
                    <RANKING order="8" place="8" resultid="12387" />
                    <RANKING order="9" place="9" resultid="12375" />
                    <RANKING order="10" place="10" resultid="12274" />
                    <RANKING order="11" place="11" resultid="12102" />
                    <RANKING order="12" place="-1" resultid="11775" />
                    <RANKING order="13" place="-1" resultid="12617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10432" agemax="54" agemin="50">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12127" />
                    <RANKING order="2" place="2" resultid="11870" />
                    <RANKING order="3" place="3" resultid="12541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10433" agemax="59" agemin="55">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10434" agemax="64" agemin="60">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="11889" />
                    <RANKING order="2" place="2" resultid="12484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10435" agemax="69" agemin="65">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12077" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10436" agemax="74" agemin="70">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12563" />
                    <RANKING order="2" place="2" resultid="12052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="10437" agemax="79" agemin="75" />
                <AGEGROUP agegroupid="10438" agemax="-1" agemin="80" />
                <AGEGROUP agegroupid="10439" agemax="-1" agemin="25">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12295" />
                    <RANKING order="2" place="2" resultid="11780" />
                    <RANKING order="3" place="3" resultid="12656" />
                    <RANKING order="4" place="4" resultid="12287" />
                    <RANKING order="5" place="5" resultid="12255" />
                    <RANKING order="6" place="6" resultid="11909" />
                    <RANKING order="7" place="7" resultid="12519" />
                    <RANKING order="8" place="8" resultid="12124" />
                    <RANKING order="9" place="9" resultid="12682" />
                    <RANKING order="10" place="10" resultid="12113" />
                    <RANKING order="11" place="11" resultid="12637" />
                    <RANKING order="12" place="12" resultid="12361" />
                    <RANKING order="13" place="13" resultid="12229" />
                    <RANKING order="14" place="14" resultid="12116" />
                    <RANKING order="15" place="15" resultid="11889" />
                    <RANKING order="16" place="16" resultid="12306" />
                    <RANKING order="17" place="17" resultid="12237" />
                    <RANKING order="18" place="18" resultid="12463" />
                    <RANKING order="19" place="19" resultid="12484" />
                    <RANKING order="20" place="20" resultid="11814" />
                    <RANKING order="21" place="21" resultid="12283" />
                    <RANKING order="22" place="22" resultid="12387" />
                    <RANKING order="23" place="23" resultid="12157" />
                    <RANKING order="24" place="24" resultid="12291" />
                    <RANKING order="25" place="25" resultid="12375" />
                    <RANKING order="26" place="26" resultid="12274" />
                    <RANKING order="27" place="27" resultid="12127" />
                    <RANKING order="28" place="28" resultid="11870" />
                    <RANKING order="29" place="29" resultid="12102" />
                    <RANKING order="30" place="30" resultid="12563" />
                    <RANKING order="31" place="31" resultid="12066" />
                    <RANKING order="32" place="32" resultid="12541" />
                    <RANKING order="33" place="33" resultid="12052" />
                    <RANKING order="34" place="34" resultid="12077" />
                    <RANKING order="35" place="-1" resultid="11775" />
                    <RANKING order="36" place="-1" resultid="12452" />
                    <RANKING order="37" place="-1" resultid="12609" />
                    <RANKING order="38" place="-1" resultid="12617" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12797" daytime="17:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12798" daytime="17:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="12799" daytime="17:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="12800" daytime="17:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="12814" daytime="17:20" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1053" daytime="17:30" gender="X" number="32" order="17" round="TIM" type="MASTERS" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="EUR" value="350" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1054" agemax="119" agemin="100" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1055" agemax="159" agemin="120" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12340" />
                    <RANKING order="2" place="2" resultid="12453" />
                    <RANKING order="3" place="-1" resultid="12410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1056" agemax="199" agemin="160" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12344" />
                    <RANKING order="2" place="2" resultid="12645" />
                    <RANKING order="3" place="3" resultid="12691" />
                    <RANKING order="4" place="4" resultid="12204" />
                    <RANKING order="5" place="5" resultid="12415" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1057" agemax="239" agemin="200" calculate="TOTAL">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="12534" />
                    <RANKING order="2" place="2" resultid="12345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1058" agemax="279" agemin="240" calculate="TOTAL" />
                <AGEGROUP agegroupid="1059" agemax="319" agemin="280" calculate="TOTAL" />
                <AGEGROUP agegroupid="1060" agemax="359" agemin="320" calculate="TOTAL" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="12801" daytime="17:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="12802" daytime="17:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="OC" nation="POR" region="ANDL" clubid="11864" name="Obidos Criativa, EEM">
          <ATHLETES>
            <ATHLETE firstname="Rui Manuel" lastname="Cunha" birthdate="1967-03-14" gender="M" nation="POR" license="210862" swrid="5418289" athleteid="11868">
              <RESULTS>
                <RESULT eventid="9737" points="264" swimtime="00:01:25.26" resultid="11869" heatid="12777" lane="7" entrytime="00:01:19.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="243" swimtime="00:00:43.86" resultid="11870" heatid="12799" lane="5" entrytime="00:00:38.63" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="José Raposo" lastname="Junior" birthdate="1963-07-27" gender="M" nation="POR" license="211457" swrid="5418281" athleteid="11871">
              <RESULTS>
                <RESULT eventid="9737" status="WDR" swimtime="00:00:00.00" resultid="11872" heatid="12777" lane="1" entrytime="00:01:20.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel Rocha" lastname="Tomás" birthdate="1983-01-27" gender="M" nation="POR" license="210528" swrid="5418282" athleteid="11873">
              <RESULTS>
                <RESULT eventid="10399" points="210" swimtime="00:00:43.17" resultid="11874" heatid="12786" lane="6" entrytime="00:00:43.56" entrycourse="LCM" />
                <RESULT eventid="9737" points="290" swimtime="00:01:17.65" resultid="11875" heatid="12777" lane="5" entrytime="00:01:19.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2203" points="236" swimtime="00:03:47.46" resultid="11876" heatid="12794" lane="1" entrytime="00:03:51.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.72" />
                    <SPLIT distance="100" swimtime="00:01:47.29" />
                    <SPLIT distance="150" swimtime="00:02:49.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo José" lastname="Amaral" birthdate="1978-10-18" gender="M" nation="POR" license="12261" swrid="4574347" athleteid="11865">
              <RESULTS>
                <RESULT eventid="9789" points="336" swimtime="00:01:31.44" resultid="11866" heatid="12790" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9737" points="375" swimtime="00:01:11.09" resultid="11867" heatid="12773" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CLIPTEAM" nation="POR" region="ANNP" clubid="11758" name="CLIP Teams Associação Desportiva" shortname="CLIP Teams">
          <ATHLETES>
            <ATHLETE firstname="Ana Monica" lastname="Eloi" birthdate="1996-12-29" gender="F" nation="POR" license="107038" swrid="4251345" athleteid="11759">
              <RESULTS>
                <RESULT eventid="2111" points="702" swimtime="00:02:33.52" resultid="11760" heatid="12736" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                    <SPLIT distance="100" swimtime="00:01:13.34" />
                    <SPLIT distance="150" swimtime="00:01:53.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1118" points="806" swimtime="00:05:22.62" resultid="11761" heatid="12769" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                    <SPLIT distance="100" swimtime="00:01:11.22" />
                    <SPLIT distance="150" swimtime="00:01:53.00" />
                    <SPLIT distance="200" swimtime="00:02:34.61" />
                    <SPLIT distance="250" swimtime="00:03:20.00" />
                    <SPLIT distance="300" swimtime="00:04:06.41" />
                    <SPLIT distance="350" swimtime="00:04:45.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2190" points="730" swimtime="00:02:50.62" resultid="11762" heatid="12792" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                    <SPLIT distance="100" swimtime="00:01:21.77" />
                    <SPLIT distance="150" swimtime="00:02:06.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10412" status="DNS" swimtime="00:00:00.00" resultid="11763" heatid="12796" lane="5" entrytime="00:00:31.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CAPGE" nation="POR" region="ANCNP" clubid="12138" name="Clube Associação de Pais da Gafanha da Encarnação" shortname="Gafanha da Encarnação">
          <ATHLETES>
            <ATHLETE firstname="Juliana Cabral" lastname="Oliveira" birthdate="1985-06-30" gender="F" nation="POR" license="131965" swrid="5045154" athleteid="12150">
              <RESULTS>
                <RESULT eventid="9605" points="294" swimtime="00:01:39.11" resultid="12151" heatid="12804" lane="1" entrytime="00:01:40.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9711" points="345" swimtime="00:01:22.34" resultid="12152" heatid="12808" lane="6" entrytime="00:01:18.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="335" swimtime="00:03:04.34" resultid="12153" heatid="12810" lane="5" entrytime="00:02:57.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                    <SPLIT distance="100" swimtime="00:01:29.04" />
                    <SPLIT distance="150" swimtime="00:02:17.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernando Duarte" lastname="Oliveira" birthdate="1986-12-19" gender="M" nation="POR" license="214457" swrid="5201379" athleteid="12146">
              <RESULTS>
                <RESULT eventid="10364" points="147" swimtime="00:00:54.64" resultid="12147" heatid="12758" lane="6" />
                <RESULT eventid="9737" points="167" swimtime="00:01:33.31" resultid="12148" heatid="12774" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9685" points="195" swimtime="00:00:39.66" resultid="12149" heatid="12743" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cristina Maria" lastname="Martins" birthdate="1971-01-03" gender="F" nation="POR" license="212345" swrid="5424167" athleteid="12142">
              <RESULTS>
                <RESULT eventid="9659" points="219" swimtime="00:00:46.93" resultid="12143" heatid="12741" lane="8" entrytime="00:00:44.75" entrycourse="SCM" />
                <RESULT eventid="10350" points="399" swimtime="00:00:48.61" resultid="12144" heatid="12757" lane="8" entrytime="00:00:50.79" entrycourse="SCM" />
                <RESULT eventid="9763" points="352" swimtime="00:01:49.15" resultid="12145" heatid="12788" lane="1" entrytime="00:01:49.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Claudio Miguel" lastname="Gomes" birthdate="1995-08-10" gender="M" nation="POR" license="105039" swrid="4251278" athleteid="12139">
              <RESULTS>
                <RESULT eventid="2177" points="699" swimtime="00:01:00.75" resultid="12140" heatid="12752" lane="4" entrytime="00:00:57.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2203" points="587" swimtime="00:02:45.27" resultid="12141" heatid="12793" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:01:19.82" />
                    <SPLIT distance="150" swimtime="00:02:03.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Manuela" lastname="Sequeira" birthdate="1968-08-13" gender="F" nation="POR" license="109962" swrid="4372593" athleteid="12158">
              <RESULTS>
                <RESULT eventid="10350" points="502" swimtime="00:00:45.04" resultid="12159" heatid="12806" lane="2" entrytime="00:00:43.70" entrycourse="LCM" />
                <RESULT eventid="9711" points="291" swimtime="00:01:31.89" resultid="12160" heatid="12808" lane="1" entrytime="00:01:29.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2190" points="494" swimtime="00:03:32.74" resultid="12161" heatid="12813" lane="4" entrytime="00:03:20.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.94" />
                    <SPLIT distance="100" swimtime="00:01:42.13" />
                    <SPLIT distance="150" swimtime="00:02:37.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rodrigo Alexandre" lastname="Ramos" birthdate="1986-04-24" gender="M" nation="BRA" license="210469" swrid="5361370" athleteid="12154">
              <RESULTS>
                <RESULT eventid="9685" points="320" swimtime="00:00:33.61" resultid="12155" heatid="12748" lane="8" entrytime="00:00:33.27" entrycourse="SCM" />
                <RESULT eventid="10364" points="223" swimtime="00:00:47.56" resultid="12156" heatid="12761" lane="1" entrytime="00:00:47.42" entrycourse="SCM" />
                <RESULT eventid="10426" points="253" swimtime="00:00:39.29" resultid="12157" heatid="12797" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="10314" swimtime="00:02:33.34" resultid="12162" heatid="12803" lane="6" entrytime="00:02:25.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.14" />
                    <SPLIT distance="100" swimtime="00:01:30.90" />
                    <SPLIT distance="150" swimtime="00:01:57.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12150" number="1" />
                    <RELAYPOSITION athleteid="12158" number="2" />
                    <RELAYPOSITION athleteid="12139" number="3" />
                    <RELAYPOSITION athleteid="12154" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="10378" swimtime="00:02:41.07" resultid="12942" heatid="12767" lane="7" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                    <SPLIT distance="100" swimtime="00:01:26.05" />
                    <SPLIT distance="150" swimtime="00:02:06.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12146" number="1" />
                    <RELAYPOSITION athleteid="12142" number="2" />
                    <RELAYPOSITION athleteid="12158" number="3" />
                    <RELAYPOSITION athleteid="12154" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SCA" nation="POR" region="ANCNP" clubid="12537" name="Sporting Clube de Aveiro">
          <ATHLETES>
            <ATHLETE firstname="Ana Maria" lastname="Martins" birthdate="1979-10-26" gender="F" nation="POR" license="123246" swrid="4756632" athleteid="12546">
              <RESULTS>
                <RESULT eventid="1144" points="250" swimtime="00:03:25.26" resultid="12547" heatid="12810" lane="6" entrytime="00:03:21.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.53" />
                    <SPLIT distance="100" swimtime="00:01:38.75" />
                    <SPLIT distance="150" swimtime="00:02:33.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9763" points="287" swimtime="00:01:54.68" resultid="12548" heatid="12787" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hugo Alexandre" lastname="Borrego" birthdate="1972-11-22" gender="M" nation="POR" license="213521" swrid="5220481" athleteid="12555">
              <RESULTS>
                <RESULT eventid="10399" status="WDR" swimtime="00:00:00.00" resultid="12556" heatid="12786" lane="1" entrytime="00:00:52.31" entrycourse="LCM" />
                <RESULT eventid="9789" status="DNS" swimtime="00:00:00.00" resultid="12557" heatid="12790" lane="6" entrytime="00:01:54.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Celso Abreu" lastname="Fernandes" birthdate="1967-11-06" gender="M" nation="POR" license="213521" swrid="5450760" athleteid="12538">
              <RESULTS>
                <RESULT eventid="9737" points="197" swimtime="00:01:34.01" resultid="12539" heatid="12775" lane="5" entrytime="00:01:41.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10399" points="176" swimtime="00:00:52.17" resultid="12540" heatid="12785" lane="4" entrytime="00:00:54.49" entrycourse="LCM" />
                <RESULT eventid="10426" points="146" swimtime="00:00:51.94" resultid="12541" heatid="12798" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jorge Vieira" lastname="Ribeiro" birthdate="1964-03-13" gender="M" nation="POR" license="128894" swrid="4939020" athleteid="12552">
              <RESULTS>
                <RESULT eventid="1157" points="415" swimtime="00:02:49.84" resultid="12553" heatid="12782" lane="6" entrytime="00:02:48.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                    <SPLIT distance="100" swimtime="00:01:23.90" />
                    <SPLIT distance="150" swimtime="00:02:07.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10399" points="254" swimtime="00:00:46.33" resultid="12554" heatid="12786" lane="5" entrytime="00:00:40.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel Castro" lastname="Trigo" birthdate="1965-11-25" gender="M" nation="POR" license="120704" swrid="4652887" athleteid="12542">
              <RESULTS>
                <RESULT eventid="9737" points="297" swimtime="00:01:26.97" resultid="12543" heatid="12777" lane="6" entrytime="00:01:23.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10399" points="186" swimtime="00:00:51.34" resultid="12544" heatid="12786" lane="7" entrytime="00:00:50.88" entrycourse="LCM" />
                <RESULT eventid="2203" points="358" swimtime="00:03:48.03" resultid="12545" heatid="12794" lane="2" entrytime="00:03:41.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.70" />
                    <SPLIT distance="100" swimtime="00:01:50.02" />
                    <SPLIT distance="150" swimtime="00:02:50.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eliana Marta" lastname="Castro" birthdate="1970-12-02" gender="F" nation="POR" license="214221" swrid="5472930" athleteid="12549">
              <RESULTS>
                <RESULT eventid="9711" points="222" swimtime="00:01:40.50" resultid="12550" heatid="12771" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10386" points="179" swimtime="00:00:55.46" resultid="12551" heatid="12784" lane="1" entrytime="00:01:01.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="10378" swimtime="00:02:40.01" resultid="12558" heatid="12767" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.38" />
                    <SPLIT distance="100" swimtime="00:01:23.51" />
                    <SPLIT distance="150" swimtime="00:02:06.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12549" number="1" />
                    <RELAYPOSITION athleteid="12538" number="2" />
                    <RELAYPOSITION athleteid="12546" number="3" />
                    <RELAYPOSITION athleteid="12552" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="CNV" nation="POR" region="ANNP" clubid="12371" name="Clube de Natacao de Valongo" shortname="Natacao de Valongo">
          <ATHLETES>
            <ATHLETE firstname="Vitor Manuel" lastname="Cardoso" birthdate="1972-12-02" gender="M" nation="POR" license="207728" swrid="4885761" athleteid="12384">
              <RESULTS>
                <RESULT eventid="9685" points="391" swimtime="00:00:32.64" resultid="12385" heatid="12748" lane="5" entrytime="00:00:31.36" entrycourse="SCM" />
                <RESULT eventid="10364" points="333" swimtime="00:00:43.69" resultid="12386" heatid="12762" lane="5" entrytime="00:00:42.33" entrycourse="SCM" />
                <RESULT eventid="10426" points="282" swimtime="00:00:39.16" resultid="12387" heatid="12799" lane="3" entrytime="00:00:40.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Paula" lastname="Santos" birthdate="1971-05-05" gender="F" nation="POR" athleteid="12403">
              <RESULTS>
                <RESULT eventid="9659" points="280" swimtime="00:00:43.23" resultid="12404" heatid="12739" lane="7" />
                <RESULT eventid="10350" points="99" swimtime="00:01:17.31" resultid="12405" heatid="12755" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Attila Janus" lastname="Ambrus" birthdate="1974-05-16" gender="M" nation="POR" license="213595" swrid="5451866" athleteid="12372">
              <RESULTS>
                <RESULT eventid="9685" points="284" swimtime="00:00:36.31" resultid="12373" heatid="12743" lane="5" />
                <RESULT eventid="9737" points="256" swimtime="00:01:23.32" resultid="12374" heatid="12774" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="243" swimtime="00:00:41.10" resultid="12375" heatid="12797" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Miguel" lastname="Ferreira" birthdate="1975-09-18" gender="M" nation="POR" license="215272" athleteid="12391">
              <RESULTS>
                <RESULT eventid="9685" status="WDR" swimtime="00:00:00.00" resultid="12392" heatid="12743" lane="3" />
                <RESULT eventid="10364" status="WDR" swimtime="00:00:00.00" resultid="12393" heatid="12759" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Filipa" lastname="Cardoso" birthdate="1992-05-07" gender="F" nation="POR" license="215209" athleteid="12380">
              <RESULTS>
                <RESULT eventid="9659" points="200" swimtime="00:00:43.24" resultid="12381" heatid="12739" lane="6" />
                <RESULT eventid="9711" points="181" swimtime="00:01:39.07" resultid="12382" heatid="12772" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10350" points="123" swimtime="00:01:03.52" resultid="12383" heatid="12755" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Susana Maria" lastname="Soares" birthdate="1970-02-19" gender="F" nation="POR" license="26158" swrid="4575644" athleteid="12406">
              <RESULTS>
                <RESULT eventid="10350" points="306" swimtime="00:00:53.11" resultid="12407" heatid="12757" lane="1" entrytime="00:00:51.45" entrycourse="LCM" />
                <RESULT eventid="9711" points="213" swimtime="00:01:42.00" resultid="12408" heatid="12772" lane="4" entrytime="00:01:42.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9763" points="308" swimtime="00:01:54.13" resultid="12409" heatid="12787" lane="4" entrytime="00:01:54.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jorge Miguel" lastname="Oliveira" birthdate="1980-05-02" gender="M" nation="POR" license="127982" swrid="4908436" athleteid="12400">
              <RESULTS>
                <RESULT eventid="9685" status="WDR" swimtime="00:00:00.00" resultid="12401" heatid="12749" lane="7" entrytime="00:00:30.66" entrycourse="SCM" />
                <RESULT eventid="1157" status="WDR" swimtime="00:00:00.00" resultid="12402" heatid="12811" lane="1" entrytime="00:02:31.23" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Joao" lastname="Mourao" birthdate="1962-12-01" gender="M" nation="POR" license="209692" swrid="5344122" athleteid="12397">
              <RESULTS>
                <RESULT eventid="9685" points="182" swimtime="00:00:45.91" resultid="12398" heatid="12745" lane="6" entrytime="00:00:44.89" entrycourse="SCM" />
                <RESULT eventid="9737" points="149" swimtime="00:01:49.23" resultid="12399" heatid="12775" lane="7" entrytime="00:01:54.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo Jorge" lastname="Fernandes" birthdate="1972-06-14" gender="M" nation="POR" license="14684" swrid="4574788" athleteid="12388">
              <RESULTS>
                <RESULT eventid="2124" points="257" swimtime="00:03:26.75" resultid="12389" heatid="12738" lane="7" entrytime="00:03:18.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.98" />
                    <SPLIT distance="100" swimtime="00:01:42.44" />
                    <SPLIT distance="150" swimtime="00:02:35.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9789" points="280" swimtime="00:01:40.95" resultid="12390" heatid="12791" lane="3" entrytime="00:01:40.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sara Gomes" lastname="Henriques" birthdate="1985-03-20" gender="F" nation="POR" license="215210" athleteid="12394">
              <RESULTS>
                <RESULT comment="609 - O(A) nadador(a) não começou a executar a viragem imediatamente após terminar a braçada na posição ventral aos 25 metros - SW 6.4" eventid="9605" status="DSQ" swimtime="00:00:00.00" resultid="12395" heatid="12733" lane="7" />
                <RESULT eventid="9659" points="217" swimtime="00:00:43.56" resultid="12396" heatid="12739" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Telmo Alexandre" lastname="Barros" birthdate="1979-12-22" gender="M" nation="POR" license="204174" swrid="4577671" athleteid="12376">
              <RESULTS>
                <RESULT eventid="9685" status="WDR" swimtime="00:00:00.00" resultid="12377" heatid="12742" lane="5" />
                <RESULT eventid="10364" status="WDR" swimtime="00:00:00.00" resultid="12378" heatid="12759" lane="6" />
                <RESULT eventid="1157" status="WDR" swimtime="00:00:00.00" resultid="12379" heatid="12780" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1053" status="WDR" swimtime="00:00:00.00" resultid="12410" heatid="12801" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12380" number="1" />
                    <RELAYPOSITION athleteid="12372" number="2" />
                    <RELAYPOSITION athleteid="12391" number="3" />
                    <RELAYPOSITION athleteid="12394" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="10378" status="WDR" swimtime="00:00:00.00" resultid="12411" heatid="12766" lane="7">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12394" number="1" />
                    <RELAYPOSITION athleteid="12384" number="2" />
                    <RELAYPOSITION athleteid="12400" number="3" />
                    <RELAYPOSITION athleteid="12380" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1061" status="WDR" swimtime="00:00:00.00" resultid="12412" heatid="12764" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12391" number="1" />
                    <RELAYPOSITION athleteid="12372" number="2" />
                    <RELAYPOSITION athleteid="12380" number="3" />
                    <RELAYPOSITION athleteid="12394" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1061" swimtime="00:06:02.34" resultid="12413" heatid="12764" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                    <SPLIT distance="100" swimtime="00:01:18.63" />
                    <SPLIT distance="150" swimtime="00:02:05.25" />
                    <SPLIT distance="200" swimtime="00:03:02.76" />
                    <SPLIT distance="250" swimtime="00:03:40.24" />
                    <SPLIT distance="300" swimtime="00:04:19.48" />
                    <SPLIT distance="350" swimtime="00:05:06.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12384" number="1" />
                    <RELAYPOSITION athleteid="12403" number="2" />
                    <RELAYPOSITION athleteid="12388" number="3" />
                    <RELAYPOSITION athleteid="12406" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="10314" swimtime="00:03:07.42" resultid="12414" heatid="12727" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                    <SPLIT distance="100" swimtime="00:01:42.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12388" number="1" />
                    <RELAYPOSITION athleteid="12380" number="2" />
                    <RELAYPOSITION athleteid="12372" number="3" />
                    <RELAYPOSITION athleteid="12394" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1053" swimtime="00:06:54.52" resultid="12415" heatid="12802" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                    <SPLIT distance="100" swimtime="00:01:34.94" />
                    <SPLIT distance="150" swimtime="00:02:29.23" />
                    <SPLIT distance="200" swimtime="00:03:32.32" />
                    <SPLIT distance="250" swimtime="00:04:17.69" />
                    <SPLIT distance="300" swimtime="00:05:12.36" />
                    <SPLIT distance="350" swimtime="00:06:02.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12388" number="1" />
                    <RELAYPOSITION athleteid="12406" number="2" />
                    <RELAYPOSITION athleteid="12384" number="3" />
                    <RELAYPOSITION athleteid="12394" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="10378" swimtime="00:02:46.81" resultid="12416" heatid="12767" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                    <SPLIT distance="100" swimtime="00:01:17.90" />
                    <SPLIT distance="150" swimtime="00:02:02.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12372" number="1" />
                    <RELAYPOSITION athleteid="12403" number="2" />
                    <RELAYPOSITION athleteid="12397" number="3" />
                    <RELAYPOSITION athleteid="12406" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="10314" swimtime="00:03:28.67" resultid="12417" heatid="12728" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.93" />
                    <SPLIT distance="100" swimtime="00:02:06.82" />
                    <SPLIT distance="150" swimtime="00:02:46.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12397" number="1" />
                    <RELAYPOSITION athleteid="12406" number="2" />
                    <RELAYPOSITION athleteid="12384" number="3" />
                    <RELAYPOSITION athleteid="12403" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="SCP" nation="POR" region="ANL" clubid="11890" name="Sporting Clube de Portugal" shortname="Sporting">
          <ATHLETES>
            <ATHLETE firstname="Paulo Paula" lastname="Carvalho" birthdate="1961-03-23" gender="M" nation="POR" license="25645" swrid="4574562" athleteid="11897">
              <RESULTS>
                <RESULT comment="Recorde Nacional " eventid="4128" points="904" swimtime="00:20:15.15" resultid="11898" heatid="12730" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                    <SPLIT distance="100" swimtime="00:01:15.17" />
                    <SPLIT distance="150" swimtime="00:01:55.38" />
                    <SPLIT distance="200" swimtime="00:02:35.97" />
                    <SPLIT distance="250" swimtime="00:03:16.79" />
                    <SPLIT distance="300" swimtime="00:03:57.71" />
                    <SPLIT distance="350" swimtime="00:04:38.70" />
                    <SPLIT distance="400" swimtime="00:05:19.70" />
                    <SPLIT distance="450" swimtime="00:06:00.47" />
                    <SPLIT distance="500" swimtime="00:06:41.03" />
                    <SPLIT distance="550" swimtime="00:07:21.64" />
                    <SPLIT distance="600" swimtime="00:08:02.32" />
                    <SPLIT distance="650" swimtime="00:08:43.40" />
                    <SPLIT distance="700" swimtime="00:09:24.30" />
                    <SPLIT distance="750" swimtime="00:10:04.93" />
                    <SPLIT distance="800" swimtime="00:10:45.30" />
                    <SPLIT distance="850" swimtime="00:11:25.85" />
                    <SPLIT distance="900" swimtime="00:12:06.54" />
                    <SPLIT distance="950" swimtime="00:12:47.14" />
                    <SPLIT distance="1000" swimtime="00:13:28.36" />
                    <SPLIT distance="1100" swimtime="00:14:50.15" />
                    <SPLIT distance="1150" swimtime="00:15:31.25" />
                    <SPLIT distance="1200" swimtime="00:16:12.04" />
                    <SPLIT distance="1250" swimtime="00:16:52.67" />
                    <SPLIT distance="1300" swimtime="00:17:34.83" />
                    <SPLIT distance="1350" swimtime="00:18:15.12" />
                    <SPLIT distance="1400" swimtime="00:18:55.44" />
                    <SPLIT distance="1450" swimtime="00:19:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Recorde Nacional " eventid="2124" points="833" swimtime="00:02:46.86" resultid="11899" heatid="12738" lane="3" entrytime="00:02:31.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:01:21.94" />
                    <SPLIT distance="150" swimtime="00:02:05.19" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="Recorde Nacional " eventid="10336" points="967" swimtime="00:02:41.51" resultid="12700" heatid="12754" lane="4" entrytime="00:02:28.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.53" />
                    <SPLIT distance="100" swimtime="00:01:16.78" />
                    <SPLIT distance="150" swimtime="00:02:00.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hugo Andre" lastname="Afonso" birthdate="1976-12-23" gender="M" nation="POR" license="204884" swrid="5216335" athleteid="11891">
              <RESULTS>
                <RESULT eventid="4128" status="WDR" swimtime="00:00:00.00" resultid="11892" />
                <RESULT eventid="9685" status="WDR" swimtime="00:00:00.00" resultid="11893" entrytime="00:00:32.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena Paula" lastname="Carvalho" birthdate="1964-05-03" gender="F" nation="POR" license="17549" swrid="4800234" athleteid="11894">
              <RESULTS>
                <RESULT eventid="4102" status="DNS" swimtime="00:00:00.00" resultid="11895" heatid="12729" lane="5" />
                <RESULT eventid="10350" points="436" swimtime="00:00:49.50" resultid="11896" heatid="12757" lane="4" entrytime="00:00:48.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CNMAIA" nation="POR" region="ANNP" clubid="12350" name="Clube de Natacao da Maia" shortname="Natacao da Maia">
          <ATHLETES>
            <ATHLETE firstname="Hugo Manuel" lastname="Ferreira" birthdate="1979-04-14" gender="M" nation="POR" athleteid="12356">
              <RESULTS>
                <RESULT eventid="1157" points="164" swimtime="00:03:26.43" resultid="12357" heatid="12780" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.03" />
                    <SPLIT distance="100" swimtime="00:01:35.03" />
                    <SPLIT distance="150" swimtime="00:02:31.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Pais" lastname="Neto" birthdate="1995-02-05" gender="M" nation="POR" license="109284" athleteid="12368">
              <RESULTS>
                <RESULT eventid="9685" points="499" swimtime="00:00:28.78" resultid="12369" heatid="12744" lane="6" />
                <RESULT eventid="9737" points="434" swimtime="00:01:04.14" resultid="12370" heatid="12774" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Pedro" lastname="Ferreira" birthdate="1995-12-25" gender="M" nation="POR" license="111411" swrid="4398286" athleteid="12358">
              <RESULTS>
                <RESULT eventid="9685" points="382" swimtime="00:00:31.47" resultid="12359" heatid="12747" lane="3" entrytime="00:00:34.04" entrycourse="SCM" />
                <RESULT eventid="10399" points="344" swimtime="00:00:35.72" resultid="12360" heatid="12786" lane="4" entrytime="00:00:36.24" entrycourse="LCM" />
                <RESULT eventid="10426" points="378" swimtime="00:00:32.75" resultid="12361" heatid="12814" lane="8" entrytime="00:00:32.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago Frederico" lastname="Dias" birthdate="1984-09-24" gender="M" nation="POR" athleteid="12354">
              <RESULTS>
                <RESULT eventid="1157" points="85" swimtime="00:04:12.81" resultid="12355" heatid="12780" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.52" />
                    <SPLIT distance="100" swimtime="00:01:55.44" />
                    <SPLIT distance="150" swimtime="00:03:04.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Pedro" lastname="Ferreira" birthdate="1964-06-30" gender="M" nation="POR" license="129087" swrid="4951641" athleteid="12362">
              <RESULTS>
                <RESULT eventid="9685" points="317" swimtime="00:00:38.15" resultid="12363" heatid="12746" lane="4" entrytime="00:00:37.91" entrycourse="LCM" />
                <RESULT eventid="10364" points="262" swimtime="00:00:47.61" resultid="12364" heatid="12761" lane="4" entrytime="00:00:45.23" entrycourse="LCM" />
                <RESULT eventid="9737" points="274" swimtime="00:01:29.27" resultid="12365" heatid="12776" lane="5" entrytime="00:01:26.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Miguel" lastname="Gomes" birthdate="1971-09-08" gender="M" nation="POR" license="214250" athleteid="12366">
              <RESULTS>
                <RESULT eventid="1157" points="346" swimtime="00:02:55.88" resultid="12367" heatid="12780" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                    <SPLIT distance="100" swimtime="00:01:24.62" />
                    <SPLIT distance="150" swimtime="00:02:12.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Pedro" lastname="Bandeira" birthdate="1995-12-20" gender="M" nation="POR" license="24291" swrid="4123339" athleteid="12351">
              <RESULTS>
                <RESULT eventid="10364" points="551" swimtime="00:00:34.46" resultid="12352" heatid="12807" lane="5" entrytime="00:00:33.85" entrycourse="LCM" />
                <RESULT eventid="9789" points="641" swimtime="00:01:11.94" resultid="12353" heatid="12790" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="GCST" nation="POR" region="ANNP" clubid="12168" name="Ginásio Clube de Santo Tirso" shortname="GCST">
          <ATHLETES>
            <ATHLETE firstname="Maria Joao" lastname="Jose" birthdate="1990-12-17" gender="F" nation="POR" license="15208" swrid="4575034" athleteid="12189">
              <RESULTS>
                <RESULT eventid="9659" points="547" swimtime="00:00:31.96" resultid="12190" heatid="12741" lane="6" entrytime="00:00:31.37" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Raquel" lastname="Lirio" birthdate="1990-12-10" gender="F" nation="POR" license="15206" swrid="4074207" athleteid="12191">
              <RESULTS>
                <RESULT eventid="1118" points="348" swimtime="00:07:04.40" resultid="12192" heatid="12769" lane="3" entrytime="00:06:59.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.84" />
                    <SPLIT distance="100" swimtime="00:01:36.10" />
                    <SPLIT distance="150" swimtime="00:02:29.80" />
                    <SPLIT distance="200" swimtime="00:03:24.95" />
                    <SPLIT distance="250" swimtime="00:04:23.68" />
                    <SPLIT distance="300" swimtime="00:05:23.67" />
                    <SPLIT distance="350" swimtime="00:06:14.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Pedro" lastname="Borges" birthdate="1974-10-31" gender="M" nation="POR" license="205247" swrid="5231495" athleteid="12179">
              <RESULTS>
                <RESULT eventid="9685" status="WDR" swimtime="00:00:00.00" resultid="12180" heatid="12742" lane="3" />
                <RESULT eventid="10364" status="WDR" swimtime="00:00:00.00" resultid="12181" heatid="12758" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Eduardo" lastname="Afonso" birthdate="1965-11-07" gender="M" nation="POR" license="207922" swrid="5032171" athleteid="12169">
              <RESULTS>
                <RESULT eventid="9685" points="306" swimtime="00:00:38.62" resultid="12170" heatid="12746" lane="3" entrytime="00:00:38.76" entrycourse="LCM" />
                <RESULT eventid="10364" points="348" swimtime="00:00:43.33" resultid="12171" heatid="12763" lane="8" entrytime="00:00:41.97" entrycourse="SCM" />
                <RESULT eventid="9789" points="336" swimtime="00:01:37.92" resultid="12172" heatid="12791" lane="5" entrytime="00:01:37.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sandra Santa" lastname="Barbara" birthdate="1975-03-22" gender="F" nation="POR" license="104504" swrid="4426885" athleteid="12176">
              <RESULTS>
                <RESULT eventid="2164" points="299" swimtime="00:01:38.74" resultid="12177" heatid="12750" lane="5" entrytime="00:01:47.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9763" points="433" swimtime="00:01:42.81" resultid="12178" heatid="12788" lane="5" entrytime="00:01:32.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cristiano Rocha" lastname="Ferreira" birthdate="1973-02-17" gender="M" nation="POR" license="131837" swrid="5041323" athleteid="12182">
              <RESULTS>
                <RESULT eventid="9685" points="260" swimtime="00:00:37.39" resultid="12183" heatid="12743" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena Manuel" lastname="Jose" birthdate="1990-12-17" gender="F" nation="POR" license="15205" swrid="4575033" athleteid="12187">
              <RESULTS>
                <RESULT eventid="9659" points="452" swimtime="00:00:34.04" resultid="12188" heatid="12741" lane="5" entrytime="00:00:30.97" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gracinda Maria" lastname="Machado" birthdate="1961-05-01" gender="F" nation="POR" license="117386" swrid="4496949" athleteid="12193">
              <RESULTS>
                <RESULT eventid="9659" points="167" swimtime="00:00:56.20" resultid="12194" heatid="12740" lane="7" entrytime="00:00:55.34" entrycourse="LCM" />
                <RESULT eventid="10386" points="171" swimtime="00:01:05.35" resultid="12195" heatid="12783" lane="5" entrytime="00:01:05.65" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariana Dias" lastname="Almeida" birthdate="1993-09-12" gender="F" nation="POR" license="22405" swrid="4074209" athleteid="12173">
              <RESULTS>
                <RESULT eventid="9659" points="534" swimtime="00:00:31.16" resultid="12174" heatid="12741" lane="4" entrytime="00:00:29.12" entrycourse="SCM" />
                <RESULT eventid="10350" points="563" swimtime="00:00:38.24" resultid="12175" heatid="12806" lane="5" entrytime="00:00:36.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno Miguel" lastname="Oliveira" birthdate="1989-05-03" gender="M" nation="POR" license="207923" swrid="5065753" athleteid="12199">
              <RESULTS>
                <RESULT eventid="9685" status="WDR" swimtime="00:00:00.00" resultid="12200" heatid="12805" lane="2" entrytime="00:00:28.43" entrycourse="LCM" />
                <RESULT eventid="9737" status="WDR" swimtime="00:00:00.00" resultid="12201" heatid="12809" lane="2" entrytime="00:01:06.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Rosario" lastname="Figueiredo" birthdate="1989-11-02" gender="M" nation="POR" license="131311" swrid="5019410" athleteid="12184">
              <RESULTS>
                <RESULT eventid="2177" points="258" swimtime="00:01:22.57" resultid="12185" heatid="12751" lane="4" entrytime="00:01:24.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="368" swimtime="00:02:28.60" resultid="12186" heatid="12811" lane="5" entrytime="00:02:22.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:11.08" />
                    <SPLIT distance="150" swimtime="00:01:50.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Augusto Mariano" lastname="Soares" birthdate="1972-03-05" gender="M" nation="POR" license="117424" swrid="4496951" athleteid="12202">
              <RESULTS>
                <RESULT comment="609 - O(A) nadador(a) não começou a executar a viragem imediatamente após terminar a braçada na posição ventral aos 25 metros - SW 6.4" eventid="2124" status="DSQ" swimtime="00:00:00.00" resultid="12203" heatid="12737" lane="5" entrytime="00:05:19.87" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Delfina Maria" lastname="Martins" birthdate="1966-11-22" gender="F" nation="POR" license="117387" swrid="4496950" athleteid="12196">
              <RESULTS>
                <RESULT eventid="9659" points="141" swimtime="00:00:55.18" resultid="12197" heatid="12740" lane="6" entrytime="00:00:52.51" entrycourse="LCM" />
                <RESULT eventid="9711" points="128" swimtime="00:02:04.26" resultid="12198" heatid="12772" lane="6" entrytime="00:01:58.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1053" swimtime="00:06:42.27" resultid="12204" heatid="12802" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.65" />
                    <SPLIT distance="100" swimtime="00:01:22.75" />
                    <SPLIT distance="150" swimtime="00:02:08.68" />
                    <SPLIT distance="200" swimtime="00:03:02.67" />
                    <SPLIT distance="250" swimtime="00:03:46.73" />
                    <SPLIT distance="300" swimtime="00:04:40.36" />
                    <SPLIT distance="350" swimtime="00:05:37.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12184" number="1" />
                    <RELAYPOSITION athleteid="12169" number="2" />
                    <RELAYPOSITION athleteid="12191" number="3" />
                    <RELAYPOSITION athleteid="12193" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="10378" status="WDR" swimtime="00:00:00.00" resultid="12205" heatid="12768" lane="4" entrytime="00:01:59.51">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12184" number="1" />
                    <RELAYPOSITION athleteid="12176" number="2" />
                    <RELAYPOSITION athleteid="12191" number="3" />
                    <RELAYPOSITION athleteid="12199" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1061" swimtime="00:05:01.71" resultid="12208" heatid="12765" lane="4" entrytime="00:04:21.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                    <SPLIT distance="100" swimtime="00:01:10.27" />
                    <SPLIT distance="150" swimtime="00:01:50.96" />
                    <SPLIT distance="200" swimtime="00:02:43.66" />
                    <SPLIT distance="250" swimtime="00:03:18.47" />
                    <SPLIT distance="300" swimtime="00:03:55.82" />
                    <SPLIT distance="350" swimtime="00:04:27.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12173" number="1" />
                    <RELAYPOSITION athleteid="12169" number="2" />
                    <RELAYPOSITION athleteid="12189" number="3" />
                    <RELAYPOSITION athleteid="12184" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="10314" swimtime="00:02:28.42" resultid="12210" heatid="12727" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.44" />
                    <SPLIT distance="100" swimtime="00:01:16.03" />
                    <SPLIT distance="150" swimtime="00:01:52.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12184" number="1" />
                    <RELAYPOSITION athleteid="12173" number="2" />
                    <RELAYPOSITION athleteid="12189" number="3" />
                    <RELAYPOSITION athleteid="12182" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="10378" swimtime="00:03:08.09" resultid="12206" heatid="12766" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="100" swimtime="00:01:34.06" />
                    <SPLIT distance="150" swimtime="00:02:12.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12169" number="1" />
                    <RELAYPOSITION athleteid="12196" number="2" />
                    <RELAYPOSITION athleteid="12182" number="3" />
                    <RELAYPOSITION athleteid="12193" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1061" status="WDR" swimtime="00:00:00.00" resultid="12207" heatid="12765" lane="7">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12169" number="1" />
                    <RELAYPOSITION athleteid="12176" number="2" />
                    <RELAYPOSITION athleteid="12179" number="3" />
                    <RELAYPOSITION athleteid="12187" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="609 - O(A) nadador(a) não começou a executar a viragem imediatamente após terminar a braçada na posição ventral aos 25 metros - SW 6.4" eventid="10314" status="DSQ" swimtime="00:00:00.00" resultid="12209" heatid="12728" lane="7">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12187" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="12179" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="12169" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="12196" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
          <COACHES>
            <COACH firstname="Sandra Santa" gender="F" lastname="Barbara" license="104504" type="HEADCOACH" />
          </COACHES>
          <OFFICIALS>
            <OFFICIAL officialid="12212" firstname="Fernando Jorge" gender="M" lastname="Vale" nation="POR" license="122112" />
          </OFFICIALS>
        </CLUB>
        <CLUB type="CLUB" code="ADP" nation="POR" region="ANNP" clubid="12418" name="Associação Desportiva de Penafiel" shortname="Penafiel">
          <ATHLETES>
            <ATHLETE firstname="Fabio Andre" lastname="Madureira" birthdate="1990-05-19" gender="M" nation="POR" license="15910" swrid="4073863" athleteid="12430">
              <RESULTS>
                <RESULT eventid="10336" points="298" swimtime="00:03:05.67" resultid="12432" heatid="12754" lane="5" entrytime="00:02:48.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                    <SPLIT distance="100" swimtime="00:01:28.80" />
                    <SPLIT distance="150" swimtime="00:02:16.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="399" swimtime="00:06:02.51" resultid="12433" heatid="12770" lane="3" entrytime="00:05:41.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:22.30" />
                    <SPLIT distance="150" swimtime="00:02:08.75" />
                    <SPLIT distance="200" swimtime="00:02:54.45" />
                    <SPLIT distance="250" swimtime="00:03:43.65" />
                    <SPLIT distance="300" swimtime="00:04:33.41" />
                    <SPLIT distance="350" swimtime="00:05:17.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9789" points="520" swimtime="00:01:16.25" resultid="12699" heatid="12812" lane="5" entrytime="00:01:12.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jaime Antonio" lastname="Soares" birthdate="1987-07-02" gender="M" nation="POR" license="208104" swrid="5320572" athleteid="12449">
              <RESULTS>
                <RESULT eventid="9632" points="213" swimtime="00:01:36.31" resultid="12450" heatid="12734" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9737" points="259" swimtime="00:01:16.90" resultid="12451" heatid="12777" lane="4" entrytime="00:01:13.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" status="WDR" swimtime="00:00:00.00" resultid="12452" heatid="12799" lane="6" entrytime="00:00:42.96" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernando Daniel" lastname="Couto" birthdate="1990-01-05" gender="M" nation="POR" license="207687" swrid="5297523" athleteid="12419">
              <RESULTS>
                <RESULT eventid="9685" status="WDR" swimtime="00:00:00.00" resultid="12420" heatid="12747" lane="4" entrytime="00:00:34.66" entrycourse="LCM" />
                <RESULT eventid="10364" status="WDR" swimtime="00:00:00.00" resultid="12421" heatid="12762" lane="6" entrytime="00:00:43.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filipe Ricardo" lastname="Dias" birthdate="1984-07-09" gender="M" nation="POR" license="207403" swrid="4005675" athleteid="12425">
              <RESULTS>
                <RESULT comment="726 - O(A) nadador(a) tocou na parede só com uma mão na chegada – SW 7.6" eventid="10364" status="DSQ" swimtime="00:00:00.00" resultid="12426" heatid="12760" lane="2" entrytime="00:00:50.43" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helder Tomas" lastname="Rocha" birthdate="1986-08-05" gender="M" nation="POR" license="203931" swrid="4235599" athleteid="12439">
              <RESULTS>
                <RESULT eventid="2177" points="208" swimtime="00:01:33.04" resultid="12440" heatid="12751" lane="5" entrytime="00:01:32.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10364" points="191" swimtime="00:00:50.10" resultid="12441" heatid="12760" lane="5" entrytime="00:00:49.69" entrycourse="SCM" />
                <RESULT eventid="1157" points="231" swimtime="00:03:01.65" resultid="12442" heatid="12782" lane="1" entrytime="00:03:04.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.87" />
                    <SPLIT distance="100" swimtime="00:01:26.55" />
                    <SPLIT distance="150" swimtime="00:02:16.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helder Daniel" lastname="Silvestre" birthdate="1980-10-20" gender="M" nation="POR" license="212657" swrid="5430596" athleteid="12446">
              <RESULTS>
                <RESULT eventid="9737" points="138" swimtime="00:01:39.13" resultid="12447" heatid="12775" lane="6" entrytime="00:01:40.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9789" points="170" swimtime="00:01:54.59" resultid="12448" heatid="12789" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Manuel" lastname="Pereira" birthdate="1972-09-01" gender="M" nation="POR" license="201104" swrid="5163399" athleteid="12436">
              <RESULTS>
                <RESULT eventid="9737" points="153" swimtime="00:01:38.83" resultid="12437" heatid="12776" lane="8" entrytime="00:01:34.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9789" points="135" swimtime="00:02:08.74" resultid="12438" heatid="12789" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anastasia" lastname="Demidova" birthdate="1993-09-27" gender="F" nation="POR" license="108673" swrid="5452924" athleteid="12422">
              <RESULTS>
                <RESULT eventid="9711" points="434" swimtime="00:01:14.07" resultid="12423" heatid="12772" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2190" points="429" swimtime="00:03:23.65" resultid="12424" heatid="12792" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.76" />
                    <SPLIT distance="100" swimtime="00:01:37.15" />
                    <SPLIT distance="150" swimtime="00:02:30.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel Paulo" lastname="Silva" birthdate="1971-05-03" gender="M" nation="POR" license="207402" swrid="4005722" athleteid="12443">
              <RESULTS>
                <RESULT eventid="9737" points="210" swimtime="00:01:32.07" resultid="12444" heatid="12776" lane="3" entrytime="00:01:30.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9789" points="261" swimtime="00:01:48.73" resultid="12445" heatid="12791" lane="7" entrytime="00:01:41.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Isabel" lastname="Ferreira" birthdate="1992-09-26" gender="F" nation="POR" license="102081" swrid="4190097" athleteid="12427">
              <RESULTS>
                <RESULT eventid="9711" points="366" swimtime="00:01:18.45" resultid="12428" heatid="12808" lane="3" entrytime="00:01:17.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2190" points="375" swimtime="00:03:33.02" resultid="12429" heatid="12813" lane="2" entrytime="00:03:34.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.83" />
                    <SPLIT distance="100" swimtime="00:01:40.34" />
                    <SPLIT distance="150" swimtime="00:02:36.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1053" swimtime="00:06:13.48" resultid="12453" heatid="12802" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.46" />
                    <SPLIT distance="100" swimtime="00:01:25.80" />
                    <SPLIT distance="150" swimtime="00:02:11.51" />
                    <SPLIT distance="200" swimtime="00:03:04.87" />
                    <SPLIT distance="250" swimtime="00:03:46.28" />
                    <SPLIT distance="300" swimtime="00:04:36.86" />
                    <SPLIT distance="350" swimtime="00:05:22.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12422" number="1" />
                    <RELAYPOSITION athleteid="12427" number="2" />
                    <RELAYPOSITION athleteid="12439" number="3" />
                    <RELAYPOSITION athleteid="12443" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="10378" swimtime="00:02:23.66" resultid="12454" heatid="12767" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:09.59" />
                    <SPLIT distance="150" swimtime="00:01:51.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12449" number="1" />
                    <RELAYPOSITION athleteid="12427" number="2" />
                    <RELAYPOSITION athleteid="12436" number="3" />
                    <RELAYPOSITION athleteid="12422" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="APUVE" nation="POR" region="ANNP" clubid="12622" name="Ass. Prop. Urbanização Vila DEste">
          <ATHLETES>
            <ATHLETE firstname="Maria Margarida" lastname="Machado" birthdate="1981-05-27" gender="F" nation="POR" license="153145" swrid="5112960" athleteid="12623">
              <RESULTS>
                <RESULT eventid="2111" points="252" swimtime="00:03:56.33" resultid="12628" heatid="12736" lane="3" entrytime="00:03:40.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.14" />
                    <SPLIT distance="100" swimtime="00:01:54.98" />
                    <SPLIT distance="150" swimtime="00:02:56.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10386" points="189" swimtime="00:00:53.18" resultid="12629" heatid="12784" lane="6" entrytime="00:00:49.22" entrycourse="SCM" />
                <RESULT eventid="1144" points="261" swimtime="00:03:22.30" resultid="12630" heatid="12810" lane="3" entrytime="00:03:13.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.75" />
                    <SPLIT distance="100" swimtime="00:01:36.41" />
                    <SPLIT distance="150" swimtime="00:02:30.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Artur Rosa" lastname="Rosa" birthdate="1976-04-01" gender="M" nation="POR" license="126945" swrid="4892368" athleteid="12625">
              <RESULTS>
                <RESULT eventid="10364" points="505" swimtime="00:00:38.02" resultid="12636" heatid="12807" lane="6" entrytime="00:00:34.09" entrycourse="SCM" />
                <RESULT eventid="10426" points="488" swimtime="00:00:32.60" resultid="12637" heatid="12814" lane="2" entrytime="00:00:30.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco Manuel" lastname="Sequeira" birthdate="1966-01-31" gender="M" nation="POR" license="201740" swrid="5180854" athleteid="12627">
              <RESULTS>
                <RESULT eventid="9632" points="198" swimtime="00:01:51.03" resultid="12638" heatid="12735" lane="7" entrytime="00:01:52.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="171" swimtime="00:03:47.89" resultid="12639" heatid="12780" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.76" />
                    <SPLIT distance="100" swimtime="00:01:45.82" />
                    <SPLIT distance="150" swimtime="00:02:46.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10364" points="317" swimtime="00:00:44.69" resultid="12640" heatid="12762" lane="8" entrytime="00:00:44.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandra Sofia" lastname="Monteiro" birthdate="1992-04-01" gender="F" nation="POR" license="15415" swrid="4269343" athleteid="12624">
              <RESULTS>
                <RESULT eventid="9605" points="595" swimtime="00:01:15.79" resultid="12631" heatid="12804" lane="4" entrytime="00:01:13.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="625" swimtime="00:02:26.22" resultid="12632" heatid="12810" lane="4" entrytime="00:02:20.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                    <SPLIT distance="100" swimtime="00:01:11.60" />
                    <SPLIT distance="150" swimtime="00:01:49.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jorge Fernando" lastname="Monteiro" birthdate="1966-02-04" gender="M" nation="POR" license="204873" athleteid="12626">
              <RESULTS>
                <RESULT eventid="9685" points="165" swimtime="00:00:47.41" resultid="12633" heatid="12743" lane="2" />
                <RESULT eventid="10364" points="77" swimtime="00:01:11.68" resultid="12634" heatid="12758" lane="1" />
                <RESULT eventid="9737" points="129" swimtime="00:01:54.62" resultid="12635" heatid="12773" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="10314" swimtime="00:02:31.18" resultid="12642" heatid="12727" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:20.65" />
                    <SPLIT distance="150" swimtime="00:01:52.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12624" number="1" />
                    <RELAYPOSITION athleteid="12627" number="2" />
                    <RELAYPOSITION athleteid="12625" number="3" />
                    <RELAYPOSITION athleteid="12623" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1061" swimtime="00:05:26.49" resultid="12643" heatid="12764" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                    <SPLIT distance="100" swimtime="00:01:05.74" />
                    <SPLIT distance="150" swimtime="00:01:47.76" />
                    <SPLIT distance="200" swimtime="00:02:34.18" />
                    <SPLIT distance="250" swimtime="00:03:22.62" />
                    <SPLIT distance="300" swimtime="00:04:20.98" />
                    <SPLIT distance="350" swimtime="00:04:52.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12624" number="1" />
                    <RELAYPOSITION athleteid="12623" number="2" />
                    <RELAYPOSITION athleteid="12627" number="3" />
                    <RELAYPOSITION athleteid="12625" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="10378" swimtime="00:02:23.45" resultid="12644" heatid="12766" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                    <SPLIT distance="100" swimtime="00:01:10.48" />
                    <SPLIT distance="150" swimtime="00:01:55.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12624" number="1" />
                    <RELAYPOSITION athleteid="12623" number="2" />
                    <RELAYPOSITION athleteid="12626" number="3" />
                    <RELAYPOSITION athleteid="12625" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1053" swimtime="00:05:52.77" resultid="12645" heatid="12802" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                    <SPLIT distance="100" swimtime="00:01:19.70" />
                    <SPLIT distance="150" swimtime="00:02:07.24" />
                    <SPLIT distance="200" swimtime="00:03:02.46" />
                    <SPLIT distance="250" swimtime="00:03:40.07" />
                    <SPLIT distance="300" swimtime="00:04:22.75" />
                    <SPLIT distance="350" swimtime="00:05:04.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12624" number="1" />
                    <RELAYPOSITION athleteid="12627" number="2" />
                    <RELAYPOSITION athleteid="12625" number="3" />
                    <RELAYPOSITION athleteid="12623" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="CDF" nation="POR" region="ANCNP" clubid="11776" name="Clube Desportivo Feirense">
          <ATHLETES>
            <ATHLETE firstname="Diana Maria" lastname="Espinheira" birthdate="1992-02-11" gender="F" nation="POR" license="103996" swrid="4123303" athleteid="11804">
              <RESULTS>
                <RESULT eventid="10350" points="405" swimtime="00:00:42.67" resultid="11805" heatid="12806" lane="7" entrytime="00:00:44.13" entrycourse="LCM" />
                <RESULT eventid="9763" points="411" swimtime="00:01:34.97" resultid="11806" heatid="12788" lane="3" entrytime="00:01:38.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filipe Jose" lastname="Baptista" birthdate="1994-01-11" gender="M" nation="POR" license="107614" swrid="4319444" athleteid="11788">
              <RESULTS>
                <RESULT eventid="9632" points="416" swimtime="00:01:13.69" resultid="11789" heatid="12734" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valdemar Silva" lastname="Paiva" birthdate="1977-09-18" gender="M" nation="POR" license="214138" swrid="5467379" athleteid="11826">
              <RESULTS>
                <RESULT eventid="9685" points="238" swimtime="00:00:37.44" resultid="11827" heatid="12746" lane="1" entrytime="00:00:40.80" entrycourse="LCM" />
                <RESULT eventid="10364" points="246" swimtime="00:00:46.35" resultid="11828" heatid="12761" lane="2" entrytime="00:00:46.81" entrycourse="LCM" />
                <RESULT eventid="9789" points="220" swimtime="00:01:45.26" resultid="11829" heatid="12791" lane="1" entrytime="00:01:45.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Lucia" lastname="Castro" birthdate="1992-12-18" gender="F" nation="POR" license="102795" swrid="4123671" athleteid="11797">
              <RESULTS>
                <RESULT eventid="10350" points="592" swimtime="00:00:37.62" resultid="11798" heatid="12806" lane="4" entrytime="00:00:36.37" entrycourse="SCM" />
                <RESULT eventid="9763" points="603" swimtime="00:01:23.62" resultid="11799" heatid="12788" lane="4" entrytime="00:01:20.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Armando Moreira" lastname="Rocha" birthdate="1974-03-19" gender="M" nation="POR" license="120744" swrid="4656165" athleteid="11830">
              <RESULTS>
                <RESULT eventid="9685" points="458" swimtime="00:00:30.96" resultid="11831" heatid="12749" lane="3" entrytime="00:00:31.02" entrycourse="LCM" />
                <RESULT eventid="10364" points="285" swimtime="00:00:46.02" resultid="11832" heatid="12762" lane="3" entrytime="00:00:43.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Paulo" lastname="Capitao" birthdate="1996-01-31" gender="M" nation="POR" license="109592" swrid="4351797" athleteid="11790">
              <RESULTS>
                <RESULT eventid="2177" points="616" swimtime="00:01:03.37" resultid="11791" heatid="12752" lane="5" entrytime="00:01:06.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10364" points="697" swimtime="00:00:31.87" resultid="11792" heatid="12759" lane="7" />
                <RESULT eventid="9789" points="607" swimtime="00:01:13.24" resultid="11793" heatid="12790" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alfredo Alexandre" lastname="Carvalho" birthdate="1973-10-24" gender="M" nation="POR" athleteid="11794">
              <RESULTS>
                <RESULT eventid="9685" points="214" swimtime="00:00:39.88" resultid="11795" heatid="12743" lane="1" />
                <RESULT eventid="9737" points="185" swimtime="00:01:32.87" resultid="11796" heatid="12774" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mario Xavier" lastname="Rocha" birthdate="1970-12-13" gender="M" nation="POR" license="202205" swrid="4135956" athleteid="11833">
              <RESULTS>
                <RESULT eventid="10364" points="350" swimtime="00:00:43.63" resultid="11834" heatid="12761" lane="5" entrytime="00:00:44.22" entrycourse="SCM" />
                <RESULT eventid="2203" points="392" swimtime="00:03:31.30" resultid="11835" heatid="12794" lane="6" entrytime="00:03:40.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.59" />
                    <SPLIT distance="100" swimtime="00:01:39.58" />
                    <SPLIT distance="150" swimtime="00:02:36.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paula Cristina" lastname="Duarte" birthdate="1965-06-02" gender="F" nation="POR" license="207732" swrid="4885556" athleteid="11800">
              <RESULTS>
                <RESULT eventid="9659" points="156" swimtime="00:00:53.30" resultid="11801" heatid="12740" lane="5" entrytime="00:00:50.15" entrycourse="SCM" />
                <RESULT eventid="10350" points="312" swimtime="00:00:55.33" resultid="11802" heatid="12756" lane="4" entrytime="00:00:52.81" entrycourse="SCM" />
                <RESULT eventid="9763" points="271" swimtime="00:02:08.46" resultid="11803" heatid="12787" lane="5" entrytime="00:01:58.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Regina Fernanda" lastname="Azevedo" birthdate="1959-11-28" gender="F" nation="POR" license="204136" swrid="5126808" athleteid="11785">
              <RESULTS>
                <RESULT eventid="9605" points="189" swimtime="00:02:21.14" resultid="11786" heatid="12733" lane="6" entrytime="00:02:17.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10350" points="155" swimtime="00:01:10.85" resultid="11787" heatid="12756" lane="6" entrytime="00:01:09.21" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Pires" lastname="Oliveira" birthdate="1969-12-21" gender="M" nation="POR" license="213336" swrid="5448810" athleteid="11817">
              <RESULTS>
                <RESULT eventid="9685" points="307" swimtime="00:00:36.62" resultid="11818" heatid="12743" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alberto Nuno" lastname="Espinheiro" birthdate="1962-08-11" gender="M" nation="POR" license="106811" swrid="4372683" athleteid="11807">
              <RESULTS>
                <RESULT eventid="9685" points="330" swimtime="00:00:37.65" resultid="11808" heatid="12747" lane="8" entrytime="00:00:36.14" entrycourse="LCM" />
                <RESULT eventid="10364" points="341" swimtime="00:00:43.64" resultid="11809" heatid="12762" lane="4" entrytime="00:00:43.24" entrycourse="LCM" />
                <RESULT eventid="9789" points="310" swimtime="00:01:40.62" resultid="11810" heatid="12791" lane="4" entrytime="00:01:37.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Paulo" lastname="Silva" birthdate="1967-02-10" gender="M" nation="POR" license="106814" swrid="4372691" athleteid="11836">
              <RESULTS>
                <RESULT eventid="9685" points="236" swimtime="00:00:39.98" resultid="11837" heatid="12746" lane="2" entrytime="00:00:39.86" entrycourse="LCM" />
                <RESULT eventid="10364" points="249" swimtime="00:00:48.84" resultid="11838" heatid="12760" lane="3" entrytime="00:00:51.05" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernando Manuel" lastname="Silva" birthdate="1969-02-28" gender="M" nation="POR" license="204631" swrid="5207456" athleteid="11839">
              <RESULTS>
                <RESULT eventid="9685" points="317" swimtime="00:00:36.25" resultid="11840" heatid="12747" lane="6" entrytime="00:00:35.45" entrycourse="LCM" />
                <RESULT eventid="10364" points="352" swimtime="00:00:43.56" resultid="11841" heatid="12763" lane="2" entrytime="00:00:41.16" entrycourse="LCM" />
                <RESULT eventid="9737" points="267" swimtime="00:01:24.94" resultid="11842" heatid="12777" lane="2" entrytime="00:01:23.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Teresa Sofia" lastname="Leite" birthdate="1992-07-31" gender="F" nation="POR" license="13596" swrid="4123273" athleteid="11815">
              <RESULTS>
                <RESULT eventid="9605" points="391" swimtime="00:01:27.17" resultid="11816" heatid="12732" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Decio Manuel" lastname="Faria" birthdate="1972-06-30" gender="M" nation="POR" license="211173" swrid="5418290" athleteid="11811">
              <RESULTS>
                <RESULT eventid="9685" points="357" swimtime="00:00:33.64" resultid="11812" heatid="12748" lane="1" entrytime="00:00:32.60" entrycourse="SCM" />
                <RESULT eventid="9789" points="332" swimtime="00:01:35.31" resultid="11813" heatid="12791" lane="6" entrytime="00:01:38.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="288" swimtime="00:00:38.87" resultid="11814" heatid="12799" lane="4" entrytime="00:00:39.32" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Liza" lastname="Orioli" birthdate="1979-06-25" gender="F" nation="POR" license="211175" swrid="5418280" athleteid="11819">
              <RESULTS>
                <RESULT eventid="9605" points="306" swimtime="00:01:40.83" resultid="11820" heatid="12804" lane="7" entrytime="00:01:44.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9763" points="388" swimtime="00:01:43.69" resultid="11821" heatid="12788" lane="7" entrytime="00:01:47.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique Silva" lastname="Paiva" birthdate="1967-04-08" gender="M" nation="POR" license="207623" swrid="5048945" athleteid="11822">
              <RESULTS>
                <RESULT eventid="9685" points="212" swimtime="00:00:41.42" resultid="11823" heatid="12745" lane="4" entrytime="00:00:42.24" entrycourse="SCM" />
                <RESULT eventid="10364" points="251" swimtime="00:00:48.71" resultid="11824" heatid="12760" lane="4" entrytime="00:00:50.38" entrycourse="LCM" />
                <RESULT eventid="9789" points="265" swimtime="00:01:48.18" resultid="11825" heatid="12790" lane="5" entrytime="00:01:50.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ruben Manuel" lastname="Almeida" birthdate="1995-08-29" gender="M" nation="POR" license="108505" swrid="4345333" athleteid="11777">
              <RESULTS>
                <RESULT eventid="10364" points="594" swimtime="00:00:33.61" resultid="11778" heatid="12807" lane="3" entrytime="00:00:34.02" entrycourse="LCM" />
                <RESULT eventid="9737" points="552" swimtime="00:00:59.21" resultid="11779" heatid="12809" lane="5" entrytime="00:01:00.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="551" swimtime="00:00:28.90" resultid="11780" heatid="12814" lane="6" entrytime="00:00:29.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="10378" swimtime="00:02:25.73" resultid="11844" heatid="12767" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:01:15.51" />
                    <SPLIT distance="150" swimtime="00:01:52.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11819" number="1" />
                    <RELAYPOSITION athleteid="11839" number="2" />
                    <RELAYPOSITION athleteid="11804" number="3" />
                    <RELAYPOSITION athleteid="11811" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT comment="Recorde Nacional " eventid="1061" swimtime="00:04:17.10" resultid="11845" heatid="12765" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.25" />
                    <SPLIT distance="100" swimtime="00:01:00.87" />
                    <SPLIT distance="150" swimtime="00:01:36.63" />
                    <SPLIT distance="200" swimtime="00:02:14.93" />
                    <SPLIT distance="250" swimtime="00:02:46.93" />
                    <SPLIT distance="300" swimtime="00:03:22.13" />
                    <SPLIT distance="350" swimtime="00:03:48.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11788" number="1" />
                    <RELAYPOSITION athleteid="11815" number="2" />
                    <RELAYPOSITION athleteid="11797" number="3" />
                    <RELAYPOSITION athleteid="11790" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="10314" swimtime="00:02:15.56" resultid="11848" heatid="12727" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:01:22.36" />
                    <SPLIT distance="150" swimtime="00:01:50.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11815" number="1" />
                    <RELAYPOSITION athleteid="11804" number="2" />
                    <RELAYPOSITION athleteid="11777" number="3" />
                    <RELAYPOSITION athleteid="11790" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="10378" swimtime="00:03:18.20" resultid="11843" heatid="12768" lane="8" entrytime="00:03:15.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.25" />
                    <SPLIT distance="100" swimtime="00:01:45.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11785" number="1" />
                    <RELAYPOSITION athleteid="11826" number="2" />
                    <RELAYPOSITION athleteid="11800" number="3" />
                    <RELAYPOSITION athleteid="11822" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="10314" swimtime="00:02:32.49" resultid="11847" heatid="12803" lane="2" entrytime="00:02:29.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.48" />
                    <SPLIT distance="100" swimtime="00:01:28.16" />
                    <SPLIT distance="150" swimtime="00:02:01.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11819" number="1" />
                    <RELAYPOSITION athleteid="11833" number="2" />
                    <RELAYPOSITION athleteid="11797" number="3" />
                    <RELAYPOSITION athleteid="11830" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="10314" swimtime="00:03:19.91" resultid="11846" heatid="12728" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.54" />
                    <SPLIT distance="100" swimtime="00:02:00.24" />
                    <SPLIT distance="150" swimtime="00:02:42.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11785" number="1" />
                    <RELAYPOSITION athleteid="11800" number="2" />
                    <RELAYPOSITION athleteid="11817" number="3" />
                    <RELAYPOSITION athleteid="11807" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="LSC" nation="POR" region="ANNP" clubid="12213" name="Leixoes Sport Club">
          <ATHLETES>
            <ATHLETE firstname="Joao Miguel" lastname="Macedo" birthdate="1974-06-03" gender="M" nation="POR" license="121593" swrid="4703142" athleteid="12279">
              <RESULTS>
                <RESULT eventid="4128" points="401" swimtime="00:22:19.55" resultid="12280" heatid="12731" lane="3" entrytime="00:21:28.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.13" />
                    <SPLIT distance="100" swimtime="00:01:18.72" />
                    <SPLIT distance="150" swimtime="00:02:02.41" />
                    <SPLIT distance="200" swimtime="00:02:46.83" />
                    <SPLIT distance="250" swimtime="00:03:31.16" />
                    <SPLIT distance="300" swimtime="00:04:15.69" />
                    <SPLIT distance="350" swimtime="00:05:00.45" />
                    <SPLIT distance="400" swimtime="00:05:45.16" />
                    <SPLIT distance="450" swimtime="00:06:29.74" />
                    <SPLIT distance="500" swimtime="00:07:14.67" />
                    <SPLIT distance="550" swimtime="00:07:59.80" />
                    <SPLIT distance="600" swimtime="00:08:44.50" />
                    <SPLIT distance="650" swimtime="00:09:29.55" />
                    <SPLIT distance="700" swimtime="00:10:15.93" />
                    <SPLIT distance="750" swimtime="00:11:01.62" />
                    <SPLIT distance="800" swimtime="00:11:46.99" />
                    <SPLIT distance="850" swimtime="00:12:32.98" />
                    <SPLIT distance="900" swimtime="00:13:18.37" />
                    <SPLIT distance="950" swimtime="00:14:04.89" />
                    <SPLIT distance="1000" swimtime="00:14:49.96" />
                    <SPLIT distance="1050" swimtime="00:15:35.12" />
                    <SPLIT distance="1100" swimtime="00:16:20.91" />
                    <SPLIT distance="1150" swimtime="00:17:06.49" />
                    <SPLIT distance="1200" swimtime="00:17:51.71" />
                    <SPLIT distance="1250" swimtime="00:18:37.16" />
                    <SPLIT distance="1300" swimtime="00:19:22.83" />
                    <SPLIT distance="1350" swimtime="00:20:08.47" />
                    <SPLIT distance="1400" swimtime="00:20:54.09" />
                    <SPLIT distance="1450" swimtime="00:21:37.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="400" swimtime="00:02:35.65" resultid="12282" heatid="12811" lane="2" entrytime="00:02:25.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                    <SPLIT distance="100" swimtime="00:01:15.35" />
                    <SPLIT distance="150" swimtime="00:01:56.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="285" swimtime="00:00:39.00" resultid="12283" heatid="12800" lane="7" entrytime="00:00:36.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filipe Monteiro" lastname="Pacheco" birthdate="1974-01-08" gender="M" nation="POR" license="130750" swrid="5003467" athleteid="12303">
              <RESULTS>
                <RESULT eventid="1157" points="379" swimtime="00:02:38.42" resultid="12304" heatid="12779" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                    <SPLIT distance="100" swimtime="00:01:14.72" />
                    <SPLIT distance="150" swimtime="00:01:56.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2203" points="454" swimtime="00:03:11.98" resultid="12305" heatid="12794" lane="5" entrytime="00:03:18.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.70" />
                    <SPLIT distance="100" swimtime="00:01:30.50" />
                    <SPLIT distance="150" swimtime="00:02:20.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="376" swimtime="00:00:35.56" resultid="12306" heatid="12798" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Luisa" lastname="Garcia" birthdate="1970-10-05" gender="F" nation="POR" license="214120" swrid="5465977" athleteid="12263">
              <RESULTS>
                <RESULT eventid="9605" points="150" swimtime="00:02:06.20" resultid="12264" heatid="12732" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10350" points="269" swimtime="00:00:55.42" resultid="12265" heatid="12756" lane="5" entrytime="00:00:54.59" entrycourse="LCM" />
                <RESULT eventid="9763" points="274" swimtime="00:01:58.68" resultid="12266" heatid="12787" lane="3" entrytime="00:02:02.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Teresa" lastname="Pinto" birthdate="1961-07-05" gender="F" nation="POR" license="120500" swrid="4638604" athleteid="12307">
              <RESULTS>
                <RESULT eventid="9605" points="245" swimtime="00:02:09.50" resultid="12308" heatid="12733" lane="3" entrytime="00:02:02.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10386" points="237" swimtime="00:00:58.63" resultid="12309" heatid="12784" lane="7" entrytime="00:00:58.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Manuela" lastname="Fonseca" birthdate="1985-05-18" gender="F" nation="POR" license="105769" swrid="4574875" athleteid="12256">
              <RESULTS>
                <RESULT eventid="9659" points="552" swimtime="00:00:31.91" resultid="12257" heatid="12739" lane="4" />
                <RESULT eventid="9711" points="498" swimtime="00:01:12.88" resultid="12258" heatid="12772" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="517" swimtime="00:02:39.60" resultid="12259" heatid="12778" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:01:17.22" />
                    <SPLIT distance="150" swimtime="00:01:58.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hugo Rafael" lastname="Guedes" birthdate="1976-10-22" gender="M" nation="POR" license="204930" swrid="5220479" athleteid="12271">
              <RESULTS>
                <RESULT eventid="9685" points="309" swimtime="00:00:35.30" resultid="12272" heatid="12747" lane="7" entrytime="00:00:35.69" entrycourse="LCM" />
                <RESULT eventid="10364" points="359" swimtime="00:00:42.60" resultid="12273" heatid="12763" lane="7" entrytime="00:00:41.93" entrycourse="LCM" />
                <RESULT eventid="10426" points="227" swimtime="00:00:42.06" resultid="12274" heatid="12798" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raquel Alexandra" lastname="Silva" birthdate="1991-06-04" gender="F" nation="POR" license="26074" swrid="4061684" athleteid="12326">
              <RESULTS>
                <RESULT eventid="1118" points="520" swimtime="00:06:11.19" resultid="12327" heatid="12769" lane="4" entrytime="00:05:58.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                    <SPLIT distance="100" swimtime="00:01:26.14" />
                    <SPLIT distance="150" swimtime="00:02:17.16" />
                    <SPLIT distance="200" swimtime="00:03:05.40" />
                    <SPLIT distance="250" swimtime="00:03:56.12" />
                    <SPLIT distance="300" swimtime="00:04:46.76" />
                    <SPLIT distance="350" swimtime="00:05:31.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10412" points="725" swimtime="00:00:31.37" resultid="12328" heatid="12796" lane="4" entrytime="00:00:30.65" entrycourse="SCM" />
                <RESULT eventid="10386" points="623" swimtime="00:00:34.91" resultid="12329" heatid="12784" lane="4" entrytime="00:00:35.56" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Manuel" lastname="Fonseca" birthdate="1987-07-18" gender="M" nation="POR" license="25159" swrid="4064552" athleteid="12252">
              <RESULTS>
                <RESULT eventid="9685" points="547" swimtime="00:00:27.05" resultid="12253" heatid="12805" lane="5" entrytime="00:00:27.55" entrycourse="LCM" />
                <RESULT eventid="9737" points="540" swimtime="00:01:00.22" resultid="12254" heatid="12773" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="474" swimtime="00:00:29.32" resultid="12255" heatid="12814" lane="7" entrytime="00:00:31.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Manuel" lastname="Baptista" birthdate="1969-09-20" gender="M" nation="POR" license="130027" swrid="4989261" athleteid="12223">
              <RESULTS>
                <RESULT eventid="10336" points="88" swimtime="00:05:11.52" resultid="12224" heatid="12754" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.56" />
                    <SPLIT distance="100" swimtime="00:02:24.94" />
                    <SPLIT distance="150" swimtime="00:03:49.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9789" points="292" swimtime="00:01:44.77" resultid="12225" heatid="12791" lane="2" entrytime="00:01:39.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2203" points="295" swimtime="00:03:52.24" resultid="12226" heatid="12794" lane="7" entrytime="00:03:45.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.40" />
                    <SPLIT distance="100" swimtime="00:01:53.22" />
                    <SPLIT distance="150" swimtime="00:02:53.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Pedro" lastname="Castro" birthdate="1974-06-10" gender="M" nation="POR" license="132355" swrid="5065798" athleteid="12234">
              <RESULTS>
                <RESULT eventid="9685" points="449" swimtime="00:00:31.15" resultid="12235" heatid="12749" lane="2" entrytime="00:00:31.72" entrycourse="LCM" />
                <RESULT eventid="9737" points="383" swimtime="00:01:12.87" resultid="12236" heatid="12809" lane="8" entrytime="00:01:12.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="335" swimtime="00:00:36.96" resultid="12237" heatid="12800" lane="2" entrytime="00:00:35.32" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Graca Maria" lastname="Almeida" birthdate="1973-08-18" gender="F" nation="POR" license="124702" swrid="4004774" athleteid="12214">
              <RESULTS>
                <RESULT eventid="9605" points="424" swimtime="00:01:30.34" resultid="12215" heatid="12804" lane="5" entrytime="00:01:28.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10412" points="483" swimtime="00:00:38.26" resultid="12216" heatid="12796" lane="3" entrytime="00:00:36.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jorge Miguel" lastname="Caselha" birthdate="1995-09-12" gender="M" nation="POR" athleteid="12230">
              <RESULTS>
                <RESULT eventid="9685" points="415" swimtime="00:00:30.62" resultid="12231" heatid="12742" lane="2" />
                <RESULT eventid="10364" points="340" swimtime="00:00:40.48" resultid="12232" heatid="12758" lane="3" />
                <RESULT eventid="9789" points="291" swimtime="00:01:33.59" resultid="12233" heatid="12789" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta Joana" lastname="Almeida" birthdate="1978-04-04" gender="F" nation="POR" athleteid="12217">
              <RESULTS>
                <RESULT eventid="10350" status="DNS" swimtime="00:00:00.00" resultid="12218" heatid="12756" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cristina Isabel" lastname="Moura" birthdate="1963-07-31" gender="F" nation="POR" license="200762" swrid="5157468" athleteid="12296">
              <RESULTS>
                <RESULT eventid="9605" points="313" swimtime="00:01:49.49" resultid="12297" heatid="12733" lane="4" entrytime="00:01:49.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10350" points="419" swimtime="00:00:50.17" resultid="12298" heatid="12757" lane="7" entrytime="00:00:50.47" entrycourse="LCM" />
                <RESULT eventid="1144" points="297" swimtime="00:03:26.36" resultid="12299" heatid="12810" lane="7" entrytime="00:03:37.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.58" />
                    <SPLIT distance="100" swimtime="00:01:37.65" />
                    <SPLIT distance="150" swimtime="00:02:32.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Bruno" lastname="Meneses" birthdate="1962-11-29" gender="M" nation="POR" license="132358" swrid="5065803" athleteid="12288">
              <RESULTS>
                <RESULT comment="611 - O(A) nadador(a) não tocou na parede com qualquer parte do corpo durante a viragem dos 75 metros - SW 6.4" eventid="9632" status="DSQ" swimtime="00:00:00.00" resultid="12289" heatid="12735" lane="5" entrytime="00:01:33.16" entrycourse="LCM" />
                <RESULT eventid="9737" points="412" swimtime="00:01:17.94" resultid="12290" heatid="12809" lane="1" entrytime="00:01:11.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="339" swimtime="00:00:40.20" resultid="12291" heatid="12800" lane="8" entrytime="00:00:36.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filipa Isabel" lastname="Reis" birthdate="1987-10-29" gender="F" nation="POR" license="153141" swrid="5112997" athleteid="12314">
              <RESULTS>
                <RESULT eventid="9659" points="240" swimtime="00:00:42.03" resultid="12315" heatid="12741" lane="1" entrytime="00:00:41.26" entrycourse="SCM" />
                <RESULT eventid="9711" points="207" swimtime="00:01:37.15" resultid="12316" heatid="12808" lane="8" entrytime="00:01:30.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10386" points="176" swimtime="00:00:53.16" resultid="12317" heatid="12784" lane="2" entrytime="00:00:51.26" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rodrigo Jorge" lastname="Rodrigues" birthdate="1969-01-20" gender="M" nation="POR" license="126944" swrid="4892367" athleteid="12318">
              <RESULTS>
                <RESULT eventid="10364" points="491" swimtime="00:00:38.98" resultid="12319" heatid="12763" lane="4" entrytime="00:00:39.47" entrycourse="LCM" />
                <RESULT eventid="9789" points="434" swimtime="00:01:31.81" resultid="12320" heatid="12812" lane="7" entrytime="00:01:27.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2203" points="400" swimtime="00:03:29.89" resultid="12321" heatid="12794" lane="3" entrytime="00:03:24.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.92" />
                    <SPLIT distance="100" swimtime="00:01:40.48" />
                    <SPLIT distance="150" swimtime="00:02:35.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sandra Marisa" lastname="Sousa" birthdate="1985-12-02" gender="F" nation="POR" license="120591" swrid="5277966" athleteid="12330">
              <RESULTS>
                <RESULT eventid="9763" points="274" swimtime="00:01:46.24" resultid="12331" heatid="12788" lane="2" entrytime="00:01:44.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10386" points="261" swimtime="00:00:48.33" resultid="12332" heatid="12784" lane="3" entrytime="00:00:48.57" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo Amorim" lastname="Rego" birthdate="1984-06-24" gender="M" nation="POR" license="15954" swrid="4064560" athleteid="12310">
              <RESULTS>
                <RESULT eventid="2124" status="WDR" swimtime="00:00:00.00" resultid="12311" heatid="12738" lane="4" entrytime="00:02:16.57" entrycourse="SCM" />
                <RESULT eventid="9685" status="WDR" swimtime="00:00:00.00" resultid="12312" heatid="12805" lane="4" entrytime="00:00:24.79" entrycourse="SCM" />
                <RESULT eventid="2177" status="WDR" swimtime="00:00:00.00" resultid="12313" heatid="12752" lane="7" entrytime="00:01:12.19" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elsa Maria" lastname="Fumega" birthdate="1978-08-21" gender="F" nation="POR" license="119665" swrid="4607079" athleteid="12260">
              <RESULTS>
                <RESULT eventid="10350" points="586" swimtime="00:00:41.03" resultid="12261" heatid="12806" lane="3" entrytime="00:00:41.85" entrycourse="LCM" />
                <RESULT eventid="10412" points="522" swimtime="00:00:36.37" resultid="12262" heatid="12796" lane="6" entrytime="00:00:36.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Antonio" lastname="Ferreira" birthdate="1958-07-17" gender="M" nation="POR" license="214085" swrid="5465976" athleteid="12248">
              <RESULTS>
                <RESULT eventid="9632" points="257" swimtime="00:01:53.48" resultid="12249" heatid="12735" lane="8" entrytime="00:02:06.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10364" points="214" swimtime="00:00:54.73" resultid="12250" heatid="12760" lane="8" entrytime="00:00:54.66" entrycourse="LCM" />
                <RESULT eventid="1157" points="283" swimtime="00:03:27.84" resultid="12251" heatid="12781" lane="3" entrytime="00:03:32.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.52" />
                    <SPLIT distance="100" swimtime="00:01:42.42" />
                    <SPLIT distance="150" swimtime="00:02:37.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Santos" lastname="Fernandes" birthdate="1962-03-28" gender="F" nation="POR" license="105263" swrid="4246947" athleteid="12242">
              <RESULTS>
                <RESULT eventid="10350" points="433" swimtime="00:00:49.61" resultid="12243" heatid="12757" lane="5" entrytime="00:00:48.96" entrycourse="LCM" />
                <RESULT eventid="1144" points="339" swimtime="00:03:17.41" resultid="12244" heatid="12778" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.65" />
                    <SPLIT distance="100" swimtime="00:01:36.12" />
                    <SPLIT distance="150" swimtime="00:02:27.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9763" points="450" swimtime="00:01:48.55" resultid="12245" heatid="12788" lane="6" entrytime="00:01:46.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nuno Duarte" lastname="Barbosa" birthdate="1996-04-07" gender="M" nation="POR" swrid="4254756" athleteid="12227">
              <RESULTS>
                <RESULT eventid="10364" points="419" swimtime="00:00:37.76" resultid="12228" heatid="12758" lane="5" />
                <RESULT eventid="10426" points="374" swimtime="00:00:32.89" resultid="12229" heatid="12797" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Miguel" lastname="Antunes" birthdate="1968-03-18" gender="M" nation="POR" license="206896" swrid="5276395" athleteid="12219">
              <RESULTS>
                <RESULT eventid="9632" points="191" swimtime="00:01:50.35" resultid="12220" heatid="12735" lane="1" entrytime="00:01:53.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2124" points="215" swimtime="00:03:51.95" resultid="12221" heatid="12737" lane="4" entrytime="00:03:49.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.11" />
                    <SPLIT distance="100" swimtime="00:01:55.17" />
                    <SPLIT distance="150" swimtime="00:02:55.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9685" points="224" swimtime="00:00:40.69" resultid="12222" heatid="12746" lane="7" entrytime="00:00:38.61" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Trigueiros" lastname="Cunha" birthdate="1964-03-27" gender="F" nation="POR" license="132357" swrid="5065800" athleteid="12238">
              <RESULTS>
                <RESULT eventid="1144" points="343" swimtime="00:03:16.71" resultid="12239" heatid="12810" lane="2" entrytime="00:03:27.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                    <SPLIT distance="100" swimtime="00:01:31.29" />
                    <SPLIT distance="150" swimtime="00:02:23.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9763" points="483" swimtime="00:01:46.06" resultid="12240" heatid="12788" lane="8" entrytime="00:01:50.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10412" points="263" swimtime="00:00:49.82" resultid="12241" heatid="12796" lane="8" entrytime="00:00:47.89" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maribel Santos" lastname="Fernandes" birthdate="1965-11-12" gender="F" nation="POR" license="26829" swrid="4574784" athleteid="12246">
              <RESULTS>
                <RESULT eventid="10350" points="509" swimtime="00:00:47.04" resultid="12247" heatid="12806" lane="1" entrytime="00:00:44.22" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernando Santos" lastname="Moreira" birthdate="1994-09-03" gender="M" nation="POR" license="15824" swrid="4561322" athleteid="12292">
              <RESULTS>
                <RESULT eventid="10336" points="443" swimtime="00:02:45.54" resultid="12293" heatid="12754" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                    <SPLIT distance="100" swimtime="00:01:14.83" />
                    <SPLIT distance="150" swimtime="00:01:58.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9737" points="532" swimtime="00:00:59.93" resultid="12294" heatid="12809" lane="4" entrytime="00:00:56.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="570" swimtime="00:00:28.58" resultid="12295" heatid="12814" lane="4" entrytime="00:00:28.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Pedro" lastname="Machado" birthdate="1986-11-09" gender="M" nation="POR" license="125910" swrid="4558986" athleteid="12284">
              <RESULTS>
                <RESULT eventid="2177" points="526" swimtime="00:01:08.37" resultid="12285" heatid="12752" lane="6" entrytime="00:01:09.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="505" swimtime="00:02:19.97" resultid="12286" heatid="12779" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                    <SPLIT distance="100" swimtime="00:01:06.42" />
                    <SPLIT distance="150" swimtime="00:01:43.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="611" swimtime="00:00:29.31" resultid="12287" heatid="12814" lane="5" entrytime="00:00:28.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Henrique" lastname="Seara" birthdate="1963-10-01" gender="M" nation="POR" license="131833" swrid="5041337" athleteid="12322">
              <RESULTS>
                <RESULT eventid="10364" points="206" swimtime="00:00:51.61" resultid="12323" heatid="12761" lane="7" entrytime="00:00:48.70" entrycourse="LCM" />
                <RESULT eventid="10399" points="123" swimtime="00:00:58.93" resultid="12324" heatid="12786" lane="8" entrytime="00:00:53.96" entrycourse="LCM" />
                <RESULT eventid="9789" points="198" swimtime="00:01:56.87" resultid="12325" heatid="12791" lane="8" entrytime="00:01:47.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anette" lastname="Kind" birthdate="1961-12-12" gender="F" nation="GER" license="120501" swrid="4648963" athleteid="12275">
              <RESULTS>
                <RESULT eventid="9711" points="248" swimtime="00:01:53.54" resultid="12276" heatid="12772" lane="5" entrytime="00:01:44.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10386" points="176" swimtime="00:01:04.70" resultid="12277" heatid="12784" lane="8" entrytime="00:01:04.22" entrycourse="SCM" />
                <RESULT eventid="2190" points="400" swimtime="00:04:14.22" resultid="12278" heatid="12813" lane="1" entrytime="00:04:11.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.89" />
                    <SPLIT distance="100" swimtime="00:02:01.73" />
                    <SPLIT distance="150" swimtime="00:03:08.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo Alexandre" lastname="Neves" birthdate="1966-04-18" gender="M" nation="POR" license="112616" swrid="4432482" athleteid="12300">
              <RESULTS>
                <RESULT eventid="4128" points="466" swimtime="00:22:41.16" resultid="12301" heatid="12731" lane="1" entrytime="00:24:20.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.54" />
                    <SPLIT distance="100" swimtime="00:01:26.82" />
                    <SPLIT distance="150" swimtime="00:02:11.86" />
                    <SPLIT distance="200" swimtime="00:02:57.10" />
                    <SPLIT distance="250" swimtime="00:03:42.62" />
                    <SPLIT distance="300" swimtime="00:04:33.89" />
                    <SPLIT distance="350" swimtime="00:05:18.25" />
                    <SPLIT distance="400" swimtime="00:06:02.97" />
                    <SPLIT distance="450" swimtime="00:06:47.55" />
                    <SPLIT distance="500" swimtime="00:07:32.33" />
                    <SPLIT distance="550" swimtime="00:08:17.26" />
                    <SPLIT distance="600" swimtime="00:09:02.02" />
                    <SPLIT distance="650" swimtime="00:09:46.68" />
                    <SPLIT distance="700" swimtime="00:10:31.92" />
                    <SPLIT distance="750" swimtime="00:11:18.11" />
                    <SPLIT distance="800" swimtime="00:12:04.30" />
                    <SPLIT distance="850" swimtime="00:12:49.65" />
                    <SPLIT distance="900" swimtime="00:13:34.84" />
                    <SPLIT distance="950" swimtime="00:14:20.51" />
                    <SPLIT distance="1000" swimtime="00:15:05.90" />
                    <SPLIT distance="1050" swimtime="00:15:50.98" />
                    <SPLIT distance="1100" swimtime="00:16:36.51" />
                    <SPLIT distance="1150" swimtime="00:17:22.21" />
                    <SPLIT distance="1200" swimtime="00:18:08.03" />
                    <SPLIT distance="1250" swimtime="00:18:53.49" />
                    <SPLIT distance="1300" swimtime="00:19:38.46" />
                    <SPLIT distance="1350" swimtime="00:20:23.88" />
                    <SPLIT distance="1400" swimtime="00:21:10.62" />
                    <SPLIT distance="1450" swimtime="00:21:57.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="412" swimtime="00:02:50.18" resultid="12302" heatid="12782" lane="3" entrytime="00:02:46.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                    <SPLIT distance="100" swimtime="00:01:22.24" />
                    <SPLIT distance="150" swimtime="00:02:06.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana DAlte" lastname="Guedes" birthdate="1980-11-23" gender="F" nation="POR" license="121739" swrid="4703108" athleteid="12267">
              <RESULTS>
                <RESULT eventid="9605" points="370" swimtime="00:01:34.66" resultid="12268" heatid="12804" lane="3" entrytime="00:01:33.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9711" points="463" swimtime="00:01:16.77" resultid="12269" heatid="12808" lane="5" entrytime="00:01:18.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10412" points="392" swimtime="00:00:40.03" resultid="12270" heatid="12796" lane="7" entrytime="00:00:38.79" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="119" agetotalmin="100" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="10378" swimtime="00:02:00.81" resultid="12333" heatid="12767" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.08" />
                    <SPLIT distance="100" swimtime="00:00:57.79" />
                    <SPLIT distance="150" swimtime="00:01:30.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12292" number="1" />
                    <RELAYPOSITION athleteid="12227" number="2" />
                    <RELAYPOSITION athleteid="12256" number="3" />
                    <RELAYPOSITION athleteid="12326" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="Recorde Nacional " eventid="1053" swimtime="00:05:24.13" resultid="12335" heatid="12801" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:01:20.47" />
                    <SPLIT distance="150" swimtime="00:02:07.10" />
                    <SPLIT distance="200" swimtime="00:03:04.74" />
                    <SPLIT distance="250" swimtime="00:03:35.25" />
                    <SPLIT distance="300" swimtime="00:04:11.57" />
                    <SPLIT distance="350" swimtime="00:04:46.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12326" number="1" />
                    <RELAYPOSITION athleteid="12330" number="2" />
                    <RELAYPOSITION athleteid="12292" number="3" />
                    <RELAYPOSITION athleteid="12230" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1061" swimtime="00:04:31.39" resultid="12334" heatid="12765" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                    <SPLIT distance="100" swimtime="00:01:01.35" />
                    <SPLIT distance="150" swimtime="00:01:37.89" />
                    <SPLIT distance="200" swimtime="00:02:18.20" />
                    <SPLIT distance="250" swimtime="00:02:52.50" />
                    <SPLIT distance="300" swimtime="00:03:30.48" />
                    <SPLIT distance="350" swimtime="00:03:59.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12284" number="1" />
                    <RELAYPOSITION athleteid="12267" number="2" />
                    <RELAYPOSITION athleteid="12256" number="3" />
                    <RELAYPOSITION athleteid="12292" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="10314" swimtime="00:02:38.07" resultid="12336" heatid="12803" lane="5" entrytime="00:02:24.30">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                    <SPLIT distance="100" swimtime="00:01:25.50" />
                    <SPLIT distance="150" swimtime="00:01:54.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12267" number="1" />
                    <RELAYPOSITION athleteid="12230" number="2" />
                    <RELAYPOSITION athleteid="12252" number="3" />
                    <RELAYPOSITION athleteid="12314" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="10314" swimtime="00:02:35.04" resultid="12337" heatid="12803" lane="3" entrytime="00:02:24.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                    <SPLIT distance="100" swimtime="00:01:25.55" />
                    <SPLIT distance="150" swimtime="00:02:04.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12214" number="1" />
                    <RELAYPOSITION athleteid="12271" number="2" />
                    <RELAYPOSITION athleteid="12260" number="3" />
                    <RELAYPOSITION athleteid="12234" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1061" swimtime="00:05:21.19" resultid="12338" heatid="12765" lane="3" entrytime="00:05:00.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                    <SPLIT distance="100" swimtime="00:01:10.90" />
                    <SPLIT distance="150" swimtime="00:01:49.31" />
                    <SPLIT distance="200" swimtime="00:02:30.73" />
                    <SPLIT distance="250" swimtime="00:03:15.23" />
                    <SPLIT distance="300" swimtime="00:04:04.88" />
                    <SPLIT distance="350" swimtime="00:04:41.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12279" number="1" />
                    <RELAYPOSITION athleteid="12260" number="2" />
                    <RELAYPOSITION athleteid="12314" number="3" />
                    <RELAYPOSITION athleteid="12318" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="10378" swimtime="00:02:09.69" resultid="12339" heatid="12768" lane="5" entrytime="00:02:07.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.95" />
                    <SPLIT distance="100" swimtime="00:01:08.00" />
                    <SPLIT distance="150" swimtime="00:01:42.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12284" number="1" />
                    <RELAYPOSITION athleteid="12314" number="2" />
                    <RELAYPOSITION athleteid="12267" number="3" />
                    <RELAYPOSITION athleteid="12252" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1053" swimtime="00:05:22.25" resultid="12340" heatid="12802" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.62" />
                    <SPLIT distance="100" swimtime="00:01:36.52" />
                    <SPLIT distance="150" swimtime="00:02:22.58" />
                    <SPLIT distance="200" swimtime="00:03:12.00" />
                    <SPLIT distance="250" swimtime="00:03:43.25" />
                    <SPLIT distance="300" swimtime="00:04:22.46" />
                    <SPLIT distance="350" swimtime="00:04:51.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12267" number="1" />
                    <RELAYPOSITION athleteid="12260" number="2" />
                    <RELAYPOSITION athleteid="12284" number="3" />
                    <RELAYPOSITION athleteid="12252" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="10378" swimtime="00:02:18.72" resultid="12341" heatid="12767" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                    <SPLIT distance="100" swimtime="00:01:07.25" />
                    <SPLIT distance="150" swimtime="00:01:43.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12234" number="1" />
                    <RELAYPOSITION athleteid="12330" number="2" />
                    <RELAYPOSITION athleteid="12260" number="3" />
                    <RELAYPOSITION athleteid="12300" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1053" swimtime="00:05:48.01" resultid="12344" heatid="12801" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.01" />
                    <SPLIT distance="100" swimtime="00:01:28.68" />
                    <SPLIT distance="150" swimtime="00:02:13.50" />
                    <SPLIT distance="200" swimtime="00:03:05.79" />
                    <SPLIT distance="250" swimtime="00:03:46.01" />
                    <SPLIT distance="300" swimtime="00:04:37.07" />
                    <SPLIT distance="350" swimtime="00:05:09.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12214" number="1" />
                    <RELAYPOSITION athleteid="12271" number="2" />
                    <RELAYPOSITION athleteid="12279" number="3" />
                    <RELAYPOSITION athleteid="12256" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1061" swimtime="00:06:05.63" resultid="12342" heatid="12764" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.26" />
                    <SPLIT distance="100" swimtime="00:01:32.56" />
                    <SPLIT distance="150" swimtime="00:02:26.56" />
                    <SPLIT distance="200" swimtime="00:03:25.82" />
                    <SPLIT distance="250" swimtime="00:04:03.85" />
                    <SPLIT distance="300" swimtime="00:04:48.61" />
                    <SPLIT distance="350" swimtime="00:05:25.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12219" number="1" />
                    <RELAYPOSITION athleteid="12263" number="2" />
                    <RELAYPOSITION athleteid="12214" number="3" />
                    <RELAYPOSITION athleteid="12300" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="10314" swimtime="00:03:19.58" resultid="12343" heatid="12728" lane="4" entrytime="00:03:11.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.81" />
                    <SPLIT distance="100" swimtime="00:01:38.23" />
                    <SPLIT distance="150" swimtime="00:02:33.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12296" number="1" />
                    <RELAYPOSITION athleteid="12246" number="2" />
                    <RELAYPOSITION athleteid="12223" number="3" />
                    <RELAYPOSITION athleteid="12322" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="1053" swimtime="00:06:46.56" resultid="12345" heatid="12802" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.09" />
                    <SPLIT distance="100" swimtime="00:01:51.39" />
                    <SPLIT distance="150" swimtime="00:02:41.73" />
                    <SPLIT distance="200" swimtime="00:03:38.75" />
                    <SPLIT distance="250" swimtime="00:04:15.77" />
                    <SPLIT distance="300" swimtime="00:04:59.59" />
                    <SPLIT distance="350" swimtime="00:05:51.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12296" number="1" />
                    <RELAYPOSITION athleteid="12238" number="2" />
                    <RELAYPOSITION athleteid="12303" number="3" />
                    <RELAYPOSITION athleteid="12322" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="10378" swimtime="00:02:43.87" resultid="12346" heatid="12768" lane="1" entrytime="00:02:36.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.86" />
                    <SPLIT distance="100" swimtime="00:01:15.64" />
                    <SPLIT distance="150" swimtime="00:02:08.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12318" number="1" />
                    <RELAYPOSITION athleteid="12223" number="2" />
                    <RELAYPOSITION athleteid="12263" number="3" />
                    <RELAYPOSITION athleteid="12214" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="4">
              <RESULTS>
                <RESULT eventid="10314" status="WDR" swimtime="00:00:00.00" resultid="12347" heatid="12803" lane="8" entrytime="00:03:08.43">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12248" number="1" />
                    <RELAYPOSITION athleteid="12242" number="2" />
                    <RELAYPOSITION athleteid="12288" number="3" />
                    <RELAYPOSITION athleteid="12307" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1061" swimtime="00:06:12.93" resultid="12348" heatid="12765" lane="2" entrytime="00:05:44.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.32" />
                    <SPLIT distance="100" swimtime="00:01:14.59" />
                    <SPLIT distance="150" swimtime="00:02:06.27" />
                    <SPLIT distance="200" swimtime="00:03:06.54" />
                    <SPLIT distance="250" swimtime="00:03:50.21" />
                    <SPLIT distance="300" swimtime="00:04:38.55" />
                    <SPLIT distance="350" swimtime="00:06:12.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12288" number="1" />
                    <RELAYPOSITION athleteid="12275" number="2" />
                    <RELAYPOSITION athleteid="12242" number="3" />
                    <RELAYPOSITION athleteid="12248" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="5">
              <RESULTS>
                <RESULT eventid="10378" swimtime="00:02:48.44" resultid="12349" heatid="12768" lane="7" entrytime="00:02:35.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:24.39" />
                    <SPLIT distance="150" swimtime="00:02:07.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12288" number="1" />
                    <RELAYPOSITION athleteid="12307" number="2" />
                    <RELAYPOSITION athleteid="12242" number="3" />
                    <RELAYPOSITION athleteid="12248" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="FCP" nation="POR" region="ANNP" clubid="12455" name="Futebol Clube do Porto" shortname="Porto">
          <ATHLETES>
            <ATHLETE firstname="Filipa Guimaraes" lastname="Goncalves" birthdate="1981-01-29" gender="F" nation="POR" athleteid="12497">
              <RESULTS>
                <RESULT eventid="9659" points="233" swimtime="00:00:44.15" resultid="12498" heatid="12739" lane="1" />
                <RESULT eventid="10350" points="194" swimtime="00:00:59.30" resultid="12499" heatid="12755" lane="3" />
                <RESULT eventid="10386" points="220" swimtime="00:00:50.59" resultid="12500" heatid="12783" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marta Prieto " lastname="Bento" birthdate="1996-02-23" gender="F" nation="POR" athleteid="12474">
              <RESULTS>
                <RESULT eventid="9659" points="254" swimtime="00:00:39.92" resultid="12475" heatid="12739" lane="3" />
                <RESULT eventid="10350" points="246" swimtime="00:00:50.38" resultid="12476" heatid="12756" lane="7" />
                <RESULT eventid="10386" points="240" swimtime="00:00:47.62" resultid="12477" heatid="12783" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo Jorge" lastname="Cohen" birthdate="1959-08-22" gender="M" nation="POR" license="26838" swrid="4319462" athleteid="12481">
              <RESULTS>
                <RESULT eventid="9685" points="572" swimtime="00:00:32.32" resultid="12482" heatid="12749" lane="1" entrytime="00:00:31.91" entrycourse="LCM" />
                <RESULT eventid="1157" points="408" swimtime="00:03:03.90" resultid="12483" heatid="12779" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.78" />
                    <SPLIT distance="150" swimtime="00:02:15.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="424" swimtime="00:00:38.78" resultid="12484" heatid="12800" lane="1" entrytime="00:00:36.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joana Azevedo Marinho Lemos" lastname="Moura" birthdate="1982-05-10" gender="F" nation="POR" license="214867" swrid="5481128" athleteid="12505">
              <RESULTS>
                <RESULT eventid="9659" points="167" swimtime="00:00:47.49" resultid="12506" heatid="12739" lane="8" />
                <RESULT comment="716 - O(A) nadador(a) não realizou  movimentos simultâneos de pernas, durante o percurso dos ... metros – SW 7.4, apos a partida" eventid="10350" status="DSQ" swimtime="00:00:00.00" resultid="12507" heatid="12755" lane="2" />
                <RESULT eventid="10386" points="134" swimtime="00:01:00.24" resultid="12508" heatid="12783" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Aderito" lastname="Chaves" birthdate="1970-10-30" gender="M" nation="POR" license="127786" swrid="4905840" athleteid="12478">
              <RESULTS>
                <RESULT eventid="2124" points="811" swimtime="00:02:29.18" resultid="12479" heatid="12738" lane="5" entrytime="00:02:26.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                    <SPLIT distance="100" swimtime="00:01:12.82" />
                    <SPLIT distance="150" swimtime="00:01:51.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="740" swimtime="00:05:32.66" resultid="12480" heatid="12770" lane="4" entrytime="00:05:32.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:12.37" />
                    <SPLIT distance="150" swimtime="00:01:56.26" />
                    <SPLIT distance="200" swimtime="00:02:39.16" />
                    <SPLIT distance="250" swimtime="00:03:28.82" />
                    <SPLIT distance="300" swimtime="00:04:16.65" />
                    <SPLIT distance="350" swimtime="00:04:55.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rosalina Bessa" lastname="Babo" birthdate="1967-02-26" gender="F" nation="POR" license="108036" swrid="4319541" athleteid="12464">
              <RESULTS>
                <RESULT eventid="10386" points="318" swimtime="00:00:45.85" resultid="12465" heatid="12784" lane="5" entrytime="00:00:44.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Jorge Leite da Silva Pei" lastname="Azevedo" birthdate="1972-06-21" gender="M" nation="POR" athleteid="12460">
              <RESULTS>
                <RESULT eventid="2177" points="258" swimtime="00:01:31.93" resultid="12461" heatid="12751" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9737" points="307" swimtime="00:01:18.40" resultid="12462" heatid="12773" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="331" swimtime="00:00:37.11" resultid="12463" heatid="12798" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cristian" lastname="Aita" birthdate="1977-11-03" gender="M" nation="POR" license="213924" swrid="5464030" athleteid="12456">
              <RESULTS>
                <RESULT eventid="4128" points="506" swimtime="00:20:51.07" resultid="12457" heatid="12730" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                    <SPLIT distance="100" swimtime="00:01:14.64" />
                    <SPLIT distance="150" swimtime="00:01:54.75" />
                    <SPLIT distance="200" swimtime="00:02:35.43" />
                    <SPLIT distance="250" swimtime="00:03:16.87" />
                    <SPLIT distance="300" swimtime="00:04:01.15" />
                    <SPLIT distance="350" swimtime="00:04:41.72" />
                    <SPLIT distance="400" swimtime="00:05:23.28" />
                    <SPLIT distance="450" swimtime="00:06:04.42" />
                    <SPLIT distance="500" swimtime="00:06:46.20" />
                    <SPLIT distance="550" swimtime="00:07:27.91" />
                    <SPLIT distance="600" swimtime="00:08:09.43" />
                    <SPLIT distance="650" swimtime="00:08:51.30" />
                    <SPLIT distance="700" swimtime="00:09:33.37" />
                    <SPLIT distance="750" swimtime="00:10:14.78" />
                    <SPLIT distance="800" swimtime="00:10:56.58" />
                    <SPLIT distance="850" swimtime="00:11:38.14" />
                    <SPLIT distance="900" swimtime="00:12:20.02" />
                    <SPLIT distance="950" swimtime="00:13:01.90" />
                    <SPLIT distance="1000" swimtime="00:13:43.85" />
                    <SPLIT distance="1050" swimtime="00:14:25.56" />
                    <SPLIT distance="1100" swimtime="00:15:07.43" />
                    <SPLIT distance="1150" swimtime="00:15:50.09" />
                    <SPLIT distance="1200" swimtime="00:16:33.07" />
                    <SPLIT distance="1250" swimtime="00:17:14.91" />
                    <SPLIT distance="1300" swimtime="00:17:56.73" />
                    <SPLIT distance="1350" swimtime="00:18:41.42" />
                    <SPLIT distance="1400" swimtime="00:19:24.05" />
                    <SPLIT distance="1450" swimtime="00:20:06.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9632" points="460" swimtime="00:01:16.46" resultid="12458" heatid="12734" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10364" points="477" swimtime="00:00:37.20" resultid="12459" heatid="12763" lane="3" entrytime="00:00:40.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia Isabel" lastname="Pereira" birthdate="1981-01-19" gender="F" nation="POR" license="106652" swrid="4507633" athleteid="12509">
              <RESULTS>
                <RESULT eventid="10350" points="482" swimtime="00:00:43.77" resultid="12510" heatid="12806" lane="6" entrytime="00:00:41.46" entrycourse="SCM" />
                <RESULT eventid="2190" points="496" swimtime="00:03:29.75" resultid="12511" heatid="12813" lane="5" entrytime="00:03:23.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.07" />
                    <SPLIT distance="100" swimtime="00:01:39.82" />
                    <SPLIT distance="150" swimtime="00:02:35.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10412" points="411" swimtime="00:00:39.38" resultid="12512" heatid="12796" lane="2" entrytime="00:00:37.01" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hugo Miguel" lastname="Vilas" birthdate="1978-11-02" gender="M" nation="POR" license="211227" swrid="4780256" athleteid="12528">
              <RESULTS>
                <RESULT eventid="9685" points="408" swimtime="00:00:31.28" resultid="12529" heatid="12749" lane="6" entrytime="00:00:31.53" entrycourse="LCM" />
                <RESULT eventid="10364" points="395" swimtime="00:00:39.61" resultid="12530" heatid="12763" lane="5" entrytime="00:00:39.65" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Alexandre" lastname="Sousa" birthdate="1982-04-09" gender="M" nation="POR" license="123374" swrid="4756745" athleteid="12524">
              <RESULTS>
                <RESULT eventid="2177" points="536" swimtime="00:01:07.94" resultid="12525" heatid="12752" lane="3" entrytime="00:01:05.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10364" points="624" swimtime="00:00:33.77" resultid="12526" heatid="12807" lane="4" entrytime="00:00:32.86" entrycourse="SCM" />
                <RESULT eventid="9789" points="617" swimtime="00:01:15.17" resultid="12527" heatid="12812" lane="4" entrytime="00:01:11.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno Miguel" lastname="Santos" birthdate="1976-07-27" gender="M" nation="POR" license="14631" swrid="4575729" athleteid="12516">
              <RESULTS>
                <RESULT eventid="1131" points="608" swimtime="00:05:41.23" resultid="12517" heatid="12770" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="150" swimtime="00:02:00.07" />
                    <SPLIT distance="200" swimtime="00:02:43.24" />
                    <SPLIT distance="250" swimtime="00:03:34.12" />
                    <SPLIT distance="300" swimtime="00:04:25.24" />
                    <SPLIT distance="350" swimtime="00:05:03.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="600" swimtime="00:02:16.01" resultid="12518" heatid="12811" lane="4" entrytime="00:02:13.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="100" swimtime="00:01:05.27" />
                    <SPLIT distance="150" swimtime="00:01:40.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="616" swimtime="00:00:30.17" resultid="12519" heatid="12814" lane="3" entrytime="00:00:29.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sandro Ricardo Costa" lastname="Ferraz" birthdate="1986-06-04" gender="M" nation="POR" athleteid="12485">
              <RESULTS>
                <RESULT eventid="9685" points="250" swimtime="00:00:36.51" resultid="12486" heatid="12743" lane="4" />
                <RESULT eventid="1157" points="185" swimtime="00:03:15.45" resultid="12487" heatid="12780" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.51" />
                    <SPLIT distance="100" swimtime="00:01:31.31" />
                    <SPLIT distance="150" swimtime="00:02:24.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9789" points="209" swimtime="00:01:47.87" resultid="12488" heatid="12789" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Manuel" lastname="Friaes" birthdate="1965-01-13" gender="F" nation="POR" license="204549" swrid="5207367" athleteid="12493">
              <RESULTS>
                <RESULT eventid="2164" points="285" swimtime="00:01:49.47" resultid="12494" heatid="12750" lane="4" entrytime="00:01:42.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10322" points="236" swimtime="00:04:17.85" resultid="12495" heatid="12753" lane="4" entrytime="00:03:56.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.66" />
                    <SPLIT distance="100" swimtime="00:02:05.05" />
                    <SPLIT distance="150" swimtime="00:03:12.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10412" points="348" swimtime="00:00:45.39" resultid="12496" heatid="12796" lane="1" entrytime="00:00:39.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vivien Patricia Ferreira" lastname="Silva" birthdate="1962-12-08" gender="F" nation="POR" license="212365" swrid="5424194" athleteid="12520">
              <RESULTS>
                <RESULT eventid="9605" points="322" swimtime="00:01:48.55" resultid="12521" heatid="12804" lane="8" entrytime="00:01:52.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9659" points="383" swimtime="00:00:39.54" resultid="12522" heatid="12740" lane="4" entrytime="00:00:45.03" entrycourse="SCM" />
                <RESULT eventid="2164" points="269" swimtime="00:01:51.66" resultid="12523" heatid="12750" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco Santos" lastname="Barros" birthdate="1972-03-17" gender="M" nation="POR" license="108661" swrid="4345381" athleteid="12466">
              <RESULTS>
                <RESULT eventid="4128" points="366" swimtime="00:23:01.82" resultid="12467" heatid="12731" lane="2" entrytime="00:23:26.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                    <SPLIT distance="100" swimtime="00:01:19.39" />
                    <SPLIT distance="150" swimtime="00:02:03.22" />
                    <SPLIT distance="200" swimtime="00:02:48.29" />
                    <SPLIT distance="250" swimtime="00:03:34.52" />
                    <SPLIT distance="300" swimtime="00:04:21.23" />
                    <SPLIT distance="350" swimtime="00:05:08.36" />
                    <SPLIT distance="400" swimtime="00:05:55.77" />
                    <SPLIT distance="450" swimtime="00:06:42.59" />
                    <SPLIT distance="500" swimtime="00:07:29.94" />
                    <SPLIT distance="550" swimtime="00:08:17.44" />
                    <SPLIT distance="600" swimtime="00:09:03.72" />
                    <SPLIT distance="650" swimtime="00:09:50.09" />
                    <SPLIT distance="700" swimtime="00:10:37.35" />
                    <SPLIT distance="750" swimtime="00:11:24.31" />
                    <SPLIT distance="800" swimtime="00:12:11.65" />
                    <SPLIT distance="850" swimtime="00:12:58.72" />
                    <SPLIT distance="900" swimtime="00:13:45.66" />
                    <SPLIT distance="950" swimtime="00:14:32.96" />
                    <SPLIT distance="1000" swimtime="00:15:20.14" />
                    <SPLIT distance="1050" swimtime="00:16:07.27" />
                    <SPLIT distance="1100" swimtime="00:16:54.41" />
                    <SPLIT distance="1150" swimtime="00:17:41.17" />
                    <SPLIT distance="1200" swimtime="00:18:27.39" />
                    <SPLIT distance="1250" swimtime="00:19:14.08" />
                    <SPLIT distance="1300" swimtime="00:20:00.15" />
                    <SPLIT distance="1350" swimtime="00:20:46.39" />
                    <SPLIT distance="1400" swimtime="00:21:32.55" />
                    <SPLIT distance="1450" swimtime="00:22:17.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9737" points="412" swimtime="00:01:11.08" resultid="12468" heatid="12809" lane="7" entrytime="00:01:10.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="363" swimtime="00:02:40.80" resultid="12469" heatid="12782" lane="4" entrytime="00:02:39.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                    <SPLIT distance="100" swimtime="00:01:17.52" />
                    <SPLIT distance="150" swimtime="00:01:59.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo Monteiro" lastname="Pinto" birthdate="1964-03-26" gender="M" nation="POR" license="211230" swrid="5425459" athleteid="12513">
              <RESULTS>
                <RESULT eventid="2124" points="114" swimtime="00:04:54.90" resultid="12514" heatid="12737" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.82" />
                    <SPLIT distance="100" swimtime="00:02:20.94" />
                    <SPLIT distance="150" swimtime="00:03:38.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="155" swimtime="00:03:55.77" resultid="12515" heatid="12781" lane="2" entrytime="00:04:04.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.22" />
                    <SPLIT distance="100" swimtime="00:01:51.28" />
                    <SPLIT distance="150" swimtime="00:02:53.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuel Filipe Martins Rocha" lastname="Ferreira" birthdate="1987-01-28" gender="M" nation="POR" athleteid="12489">
              <RESULTS>
                <RESULT eventid="9685" points="312" swimtime="00:00:32.61" resultid="12490" heatid="12744" lane="1" />
                <RESULT eventid="10364" points="219" swimtime="00:00:46.13" resultid="12491" heatid="12759" lane="2" />
                <RESULT eventid="9737" points="272" swimtime="00:01:15.67" resultid="12492" heatid="12775" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mario Jorge" lastname="Barros" birthdate="1956-06-06" gender="M" nation="POR" license="128252" swrid="4913068" athleteid="12470">
              <RESULTS>
                <RESULT eventid="9632" points="334" swimtime="00:01:44.29" resultid="12471" heatid="12735" lane="6" entrytime="00:01:45.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10364" points="470" swimtime="00:00:43.65" resultid="12472" heatid="12762" lane="7" entrytime="00:00:43.09" entrycourse="SCM" />
                <RESULT comment="609 - O(A) nadador(a) não começou a executar a viragem imediatamente após terminar a braçada na posição ventral aos 25 metros - SW 6.4" eventid="10399" status="DSQ" swimtime="00:00:00.00" resultid="12473" heatid="12785" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alfredo Coelho" lastname="Magalhaes" birthdate="1953-11-29" gender="M" nation="POR" license="210499" swrid="5365300" athleteid="12501">
              <RESULTS>
                <RESULT eventid="9685" points="87" swimtime="00:01:02.23" resultid="12502" heatid="12744" lane="3" entrytime="00:01:03.78" entrycourse="SCM" />
                <RESULT eventid="9737" points="88" swimtime="00:02:17.27" resultid="12503" heatid="12775" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.56" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="723 - O(A) nadador(a) tocou só com uma mão na parede na viragem dos 25 metros – SW 7.6" eventid="2203" status="DSQ" swimtime="00:00:00.00" resultid="12504" heatid="12793" lane="6" entrytime="00:04:45.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="10378" swimtime="00:02:19.88" resultid="12531" heatid="12766" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                    <SPLIT distance="100" swimtime="00:01:06.23" />
                    <SPLIT distance="150" swimtime="00:01:45.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12466" number="1" />
                    <RELAYPOSITION athleteid="12489" number="2" />
                    <RELAYPOSITION athleteid="12474" number="3" />
                    <RELAYPOSITION athleteid="12509" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="1061" swimtime="00:05:02.19" resultid="12532" heatid="12764" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                    <SPLIT distance="100" swimtime="00:01:03.51" />
                    <SPLIT distance="150" swimtime="00:01:40.58" />
                    <SPLIT distance="200" swimtime="00:02:23.31" />
                    <SPLIT distance="250" swimtime="00:02:55.04" />
                    <SPLIT distance="300" swimtime="00:03:28.82" />
                    <SPLIT distance="350" swimtime="00:04:13.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12524" number="1" />
                    <RELAYPOSITION athleteid="12509" number="2" />
                    <RELAYPOSITION athleteid="12478" number="3" />
                    <RELAYPOSITION athleteid="12493" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="10314" swimtime="00:03:04.58" resultid="12533" heatid="12728" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.60" />
                    <SPLIT distance="100" swimtime="00:01:38.02" />
                    <SPLIT distance="150" swimtime="00:02:16.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12497" number="1" />
                    <RELAYPOSITION athleteid="12485" number="2" />
                    <RELAYPOSITION athleteid="12460" number="3" />
                    <RELAYPOSITION athleteid="12505" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="4">
              <RESULTS>
                <RESULT comment="Recorde Nacional " eventid="1053" swimtime="00:05:45.20" resultid="12534" heatid="12802" lane="4" entrytime="00:05:30.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                    <SPLIT distance="100" swimtime="00:01:08.91" />
                    <SPLIT distance="150" swimtime="00:01:43.49" />
                    <SPLIT distance="200" swimtime="00:02:21.69" />
                    <SPLIT distance="250" swimtime="00:03:12.06" />
                    <SPLIT distance="350" swimtime="00:04:55.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12478" number="1" />
                    <RELAYPOSITION athleteid="12524" number="2" />
                    <RELAYPOSITION athleteid="12493" number="3" />
                    <RELAYPOSITION athleteid="12520" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="279" agetotalmin="240" gender="X" number="5">
              <RESULTS>
                <RESULT eventid="10378" swimtime="00:02:30.70" resultid="12535" heatid="12768" lane="3" entrytime="00:02:26.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="100" swimtime="00:01:11.85" />
                    <SPLIT distance="150" swimtime="00:01:50.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12481" number="1" />
                    <RELAYPOSITION athleteid="12493" number="2" />
                    <RELAYPOSITION athleteid="12470" number="3" />
                    <RELAYPOSITION athleteid="12520" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="10314" swimtime="00:03:14.64" resultid="12536" heatid="12803" lane="1" entrytime="00:02:55.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.80" />
                    <SPLIT distance="100" swimtime="00:01:50.51" />
                    <SPLIT distance="150" swimtime="00:02:39.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12493" number="1" />
                    <RELAYPOSITION athleteid="12501" number="2" />
                    <RELAYPOSITION athleteid="12520" number="3" />
                    <RELAYPOSITION athleteid="12481" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="GDNFAMA" nation="POR" region="ANNP" clubid="11960" name="Grupo Desportivo Natação de V.N.Famalicão" shortname="Famalicão">
          <ATHLETES>
            <ATHLETE firstname="Antonio Sergio" lastname="Costa" birthdate="1984-03-23" gender="M" nation="POR" license="214235" swrid="4564417" athleteid="12649">
              <RESULTS>
                <RESULT eventid="10364" points="582" swimtime="00:00:34.57" resultid="12650" heatid="12807" lane="1" entrytime="00:00:36.79" entrycourse="LCM" />
                <RESULT eventid="9789" points="595" swimtime="00:01:16.08" resultid="12651" heatid="12812" lane="6" entrytime="00:01:22.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2203" points="520" swimtime="00:02:54.80" resultid="12652" heatid="12794" lane="4" entrytime="00:03:09.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                    <SPLIT distance="100" swimtime="00:01:21.54" />
                    <SPLIT distance="150" swimtime="00:02:07.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisca Silva" lastname="Carmo" birthdate="1994-09-20" gender="F" nation="POR" license="15615" swrid="4574532" athleteid="12646">
              <RESULTS>
                <RESULT eventid="9605" points="425" swimtime="00:01:24.78" resultid="12647" heatid="12732" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10386" points="415" swimtime="00:00:39.69" resultid="12648" heatid="12783" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cristina Alexandra" lastname="Furtado" birthdate="1996-02-22" gender="F" nation="POR" license="110596" swrid="4375304" athleteid="12657">
              <RESULTS>
                <RESULT eventid="9659" points="561" swimtime="00:00:30.65" resultid="12658" heatid="12739" lane="5" />
                <RESULT eventid="9711" points="545" swimtime="00:01:08.68" resultid="12659" heatid="12771" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10412" points="463" swimtime="00:00:35.93" resultid="12660" heatid="12795" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luís Manuel" lastname="Oliveira" birthdate="1988-12-02" gender="M" nation="POR" license="215275" athleteid="12665">
              <RESULTS>
                <RESULT eventid="9685" points="395" swimtime="00:00:30.14" resultid="12666" heatid="12744" lane="7" />
                <RESULT eventid="10364" points="427" swimtime="00:00:36.93" resultid="12667" heatid="12758" lane="8" />
                <RESULT eventid="9737" points="354" swimtime="00:01:09.26" resultid="12668" heatid="12774" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco Zamith" lastname="Passos" birthdate="1983-12-21" gender="M" nation="POR" license="18082" swrid="4564418" athleteid="12669">
              <RESULTS>
                <RESULT eventid="2177" points="573" swimtime="00:01:06.45" resultid="12670" heatid="12751" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="628" swimtime="00:02:10.16" resultid="12672" heatid="12781" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                    <SPLIT distance="100" swimtime="00:01:02.49" />
                    <SPLIT distance="150" swimtime="00:01:36.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4128" points="628" swimtime="00:19:29.68" resultid="12673" heatid="12730" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="100" swimtime="00:01:07.66" />
                    <SPLIT distance="150" swimtime="00:01:45.06" />
                    <SPLIT distance="200" swimtime="00:02:22.93" />
                    <SPLIT distance="250" swimtime="00:03:00.90" />
                    <SPLIT distance="300" swimtime="00:03:39.49" />
                    <SPLIT distance="350" swimtime="00:04:17.79" />
                    <SPLIT distance="400" swimtime="00:04:56.60" />
                    <SPLIT distance="450" swimtime="00:05:35.65" />
                    <SPLIT distance="500" swimtime="00:06:15.23" />
                    <SPLIT distance="550" swimtime="00:06:54.55" />
                    <SPLIT distance="600" swimtime="00:07:34.14" />
                    <SPLIT distance="650" swimtime="00:08:13.90" />
                    <SPLIT distance="700" swimtime="00:08:54.26" />
                    <SPLIT distance="750" swimtime="00:09:34.03" />
                    <SPLIT distance="800" swimtime="00:10:13.86" />
                    <SPLIT distance="850" swimtime="00:10:53.53" />
                    <SPLIT distance="900" swimtime="00:11:33.56" />
                    <SPLIT distance="950" swimtime="00:12:13.40" />
                    <SPLIT distance="1000" swimtime="00:12:53.10" />
                    <SPLIT distance="1050" swimtime="00:13:33.16" />
                    <SPLIT distance="1100" swimtime="00:14:12.73" />
                    <SPLIT distance="1150" swimtime="00:14:52.10" />
                    <SPLIT distance="1200" swimtime="00:15:32.54" />
                    <SPLIT distance="1250" swimtime="00:16:12.61" />
                    <SPLIT distance="1300" swimtime="00:16:52.92" />
                    <SPLIT distance="1350" swimtime="00:17:32.40" />
                    <SPLIT distance="1400" swimtime="00:18:12.18" />
                    <SPLIT distance="1450" swimtime="00:18:52.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mario Rui" lastname="Cunha" birthdate="1993-01-06" gender="M" nation="POR" license="15611" swrid="4574699" athleteid="12653">
              <RESULTS>
                <RESULT eventid="9685" points="568" swimtime="00:00:27.57" resultid="12654" heatid="12742" lane="6" />
                <RESULT eventid="9737" points="456" swimtime="00:01:03.08" resultid="12655" heatid="12774" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="535" swimtime="00:00:29.18" resultid="12656" heatid="12798" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nuno Miguel" lastname="Macedo" birthdate="1982-06-29" gender="M" nation="POR" license="23308" swrid="4061678" athleteid="12661">
              <RESULTS>
                <RESULT eventid="9685" points="503" swimtime="00:00:28.92" resultid="12662" heatid="12805" lane="7" entrytime="00:00:28.70" entrycourse="LCM" />
                <RESULT eventid="9737" points="480" swimtime="00:01:05.65" resultid="12663" heatid="12809" lane="3" entrytime="00:01:05.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10364" points="562" swimtime="00:00:34.97" resultid="12664" heatid="12807" lane="2" entrytime="00:00:35.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="10314" swimtime="00:02:13.30" resultid="11989" heatid="12728" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:14.23" />
                    <SPLIT distance="150" swimtime="00:01:42.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12646" number="1" />
                    <RELAYPOSITION athleteid="12649" number="2" />
                    <RELAYPOSITION athleteid="12669" number="3" />
                    <RELAYPOSITION athleteid="12657" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="10378" swimtime="00:02:03.00" resultid="11990" heatid="12766" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                    <SPLIT distance="100" swimtime="00:01:03.03" />
                    <SPLIT distance="150" swimtime="00:01:32.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12661" number="1" />
                    <RELAYPOSITION athleteid="12646" number="2" />
                    <RELAYPOSITION athleteid="12665" number="3" />
                    <RELAYPOSITION athleteid="12657" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="CFV" nation="POR" region="ANNP" clubid="11905" name="Clube Fluvial Vilacondense" shortname="Vilacondense">
          <ATHLETES>
            <ATHLETE firstname="Joaquim Silva" lastname="Santos" birthdate="1965-09-01" gender="M" nation="POR" license="153262" swrid="5115804" athleteid="12687">
              <RESULTS>
                <RESULT comment="603 - O(A) nadador(a) abandonou a posição dorsal durante o percurso dos 45 metros – SW 6.2" eventid="10399" status="DSQ" swimtime="00:00:00.00" resultid="12688" heatid="12785" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno Santos" lastname="Maia" birthdate="1981-08-09" gender="M" nation="POR" license="212423" swrid="5424166" athleteid="12679">
              <RESULTS>
                <RESULT eventid="2177" points="482" swimtime="00:01:12.18" resultid="12680" heatid="12752" lane="1" entrytime="00:01:12.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" status="DNS" swimtime="00:00:00.00" resultid="12681" heatid="12811" lane="6" entrytime="00:02:23.40" entrycourse="SCM" />
                <RESULT eventid="10426" points="532" swimtime="00:00:31.01" resultid="12682" heatid="12814" lane="1" entrytime="00:00:31.06" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Maria" lastname="Soares" birthdate="1971-01-14" gender="F" nation="POR" license="153261" swrid="5115809" athleteid="12689">
              <RESULTS>
                <RESULT eventid="10386" points="94" swimtime="00:01:08.61" resultid="12690" heatid="12783" lane="4" entrytime="00:01:05.22" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Renato Pereira" lastname="Neiva" birthdate="1989-11-12" gender="M" nation="POR" license="104826" athleteid="11913">
              <RESULTS>
                <RESULT eventid="4128" points="359" swimtime="00:23:00.80" resultid="11914" heatid="12730" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:11.92" />
                    <SPLIT distance="150" swimtime="00:01:55.03" />
                    <SPLIT distance="200" swimtime="00:02:38.76" />
                    <SPLIT distance="250" swimtime="00:03:23.80" />
                    <SPLIT distance="300" swimtime="00:04:09.54" />
                    <SPLIT distance="350" swimtime="00:04:56.32" />
                    <SPLIT distance="400" swimtime="00:05:43.32" />
                    <SPLIT distance="450" swimtime="00:06:29.95" />
                    <SPLIT distance="500" swimtime="00:07:16.35" />
                    <SPLIT distance="550" swimtime="00:08:02.89" />
                    <SPLIT distance="600" swimtime="00:08:49.56" />
                    <SPLIT distance="650" swimtime="00:09:36.94" />
                    <SPLIT distance="700" swimtime="00:10:23.43" />
                    <SPLIT distance="750" swimtime="00:11:10.32" />
                    <SPLIT distance="800" swimtime="00:11:58.06" />
                    <SPLIT distance="850" swimtime="00:12:45.54" />
                    <SPLIT distance="900" swimtime="00:13:32.38" />
                    <SPLIT distance="950" swimtime="00:14:20.36" />
                    <SPLIT distance="1000" swimtime="00:15:07.63" />
                    <SPLIT distance="1050" swimtime="00:15:55.70" />
                    <SPLIT distance="1100" swimtime="00:16:43.67" />
                    <SPLIT distance="1150" swimtime="00:17:32.51" />
                    <SPLIT distance="1200" swimtime="00:18:21.16" />
                    <SPLIT distance="1250" swimtime="00:19:09.12" />
                    <SPLIT distance="1300" swimtime="00:19:55.85" />
                    <SPLIT distance="1350" swimtime="00:20:42.76" />
                    <SPLIT distance="1400" swimtime="00:21:29.50" />
                    <SPLIT distance="1450" swimtime="00:22:16.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10364" points="373" swimtime="00:00:38.62" resultid="11915" heatid="12758" lane="2" />
                <RESULT eventid="1157" points="321" swimtime="00:02:35.44" resultid="11916" heatid="12780" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="100" swimtime="00:01:13.09" />
                    <SPLIT distance="150" swimtime="00:01:55.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Catarina Teixeira" lastname="Esteves" birthdate="1978-01-26" gender="F" nation="POR" license="111258" athleteid="12676">
              <RESULTS>
                <RESULT eventid="9711" points="544" swimtime="00:01:12.77" resultid="12677" heatid="12771" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9763" points="459" swimtime="00:01:38.10" resultid="12678" heatid="12787" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago Dourado" lastname="Campos" birthdate="1988-09-06" gender="M" nation="POR" license="23051" swrid="4064368" athleteid="11906">
              <RESULTS>
                <RESULT eventid="9685" points="542" swimtime="00:00:27.13" resultid="11907" heatid="12742" lane="7" />
                <RESULT eventid="9737" points="477" swimtime="00:01:02.74" resultid="11908" heatid="12774" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="438" swimtime="00:00:30.11" resultid="11909" heatid="12797" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Debora Filipa" lastname="Santos" birthdate="1992-06-17" gender="F" nation="POR" license="132091" swrid="5098198" athleteid="12683">
              <RESULTS>
                <RESULT eventid="9659" points="73" swimtime="00:01:00.34" resultid="12684" heatid="12740" lane="1" entrytime="00:01:00.00" entrycourse="SCM" />
                <RESULT eventid="1144" points="99" swimtime="00:04:30.12" resultid="12685" heatid="12778" lane="4" entrytime="00:04:27.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.32" />
                    <SPLIT distance="100" swimtime="00:02:12.15" />
                    <SPLIT distance="150" swimtime="00:03:22.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10412" points="30" swimtime="00:01:29.30" resultid="12686" heatid="12795" lane="3" entrytime="00:01:20.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1053" swimtime="00:06:12.30" resultid="12691" heatid="12802" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.44" />
                    <SPLIT distance="100" swimtime="00:01:28.98" />
                    <SPLIT distance="150" swimtime="00:02:08.88" />
                    <SPLIT distance="200" swimtime="00:02:57.37" />
                    <SPLIT distance="250" swimtime="00:03:31.66" />
                    <SPLIT distance="300" swimtime="00:04:10.36" />
                    <SPLIT distance="350" swimtime="00:05:05.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12676" number="1" />
                    <RELAYPOSITION athleteid="11913" number="2" />
                    <RELAYPOSITION athleteid="12679" number="3" />
                    <RELAYPOSITION athleteid="12689" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="10378" swimtime="00:02:24.89" resultid="12692" heatid="12766" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                    <SPLIT distance="100" swimtime="00:01:00.64" />
                    <SPLIT distance="150" swimtime="00:01:32.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12679" number="1" />
                    <RELAYPOSITION athleteid="11913" number="2" />
                    <RELAYPOSITION athleteid="12676" number="3" />
                    <RELAYPOSITION athleteid="12689" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="UDO" nation="POR" region="ANCNP" clubid="12584" name="UD Oliveirense/FERSILVA" />
        <CLUB type="CLUB" code="SAD" nation="POR" region="ANL" clubid="11885" name="Sport Algés e Dafundo">
          <ATHLETES>
            <ATHLETE firstname="Jaime Carlos" lastname="Bento" birthdate="1961-03-05" gender="M" nation="POR" license="118614" swrid="4583590" athleteid="11886">
              <RESULTS>
                <RESULT eventid="4128" points="860" swimtime="00:20:35.47" resultid="11887" heatid="12730" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:15.80" />
                    <SPLIT distance="150" swimtime="00:01:56.52" />
                    <SPLIT distance="200" swimtime="00:02:37.59" />
                    <SPLIT distance="250" swimtime="00:03:18.79" />
                    <SPLIT distance="300" swimtime="00:04:00.05" />
                    <SPLIT distance="350" swimtime="00:04:41.70" />
                    <SPLIT distance="400" swimtime="00:05:23.45" />
                    <SPLIT distance="450" swimtime="00:06:05.00" />
                    <SPLIT distance="500" swimtime="00:06:46.28" />
                    <SPLIT distance="550" swimtime="00:07:27.93" />
                    <SPLIT distance="600" swimtime="00:08:09.67" />
                    <SPLIT distance="650" swimtime="00:08:51.18" />
                    <SPLIT distance="700" swimtime="00:09:32.74" />
                    <SPLIT distance="750" swimtime="00:10:14.31" />
                    <SPLIT distance="800" swimtime="00:10:55.85" />
                    <SPLIT distance="850" swimtime="00:11:37.28" />
                    <SPLIT distance="900" swimtime="00:12:19.12" />
                    <SPLIT distance="950" swimtime="00:13:00.52" />
                    <SPLIT distance="1000" swimtime="00:13:42.30" />
                    <SPLIT distance="1050" swimtime="00:14:23.81" />
                    <SPLIT distance="1100" swimtime="00:15:06.20" />
                    <SPLIT distance="1150" swimtime="00:15:47.98" />
                    <SPLIT distance="1200" swimtime="00:16:30.17" />
                    <SPLIT distance="1250" swimtime="00:17:11.48" />
                    <SPLIT distance="1300" swimtime="00:17:53.53" />
                    <SPLIT distance="1350" swimtime="00:18:34.85" />
                    <SPLIT distance="1400" swimtime="00:19:16.09" />
                    <SPLIT distance="1450" swimtime="00:19:57.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="797" swimtime="00:02:27.17" resultid="11888" heatid="12811" lane="7" entrytime="00:02:30.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                    <SPLIT distance="100" swimtime="00:01:10.81" />
                    <SPLIT distance="150" swimtime="00:01:49.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="573" swimtime="00:00:35.09" resultid="11889" heatid="12800" lane="6" entrytime="00:00:34.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CGA" nation="POR" region="ANCNP" clubid="12163" name="Clube dos Galitos / Bresimar" shortname="Galitos / Bresimar">
          <ATHLETES>
            <ATHLETE firstname="Joana Isabel" lastname="Cunha" birthdate="1980-07-17" gender="F" nation="POR" license="117125" swrid="4475974" athleteid="12164">
              <RESULTS>
                <RESULT eventid="9659" points="620" swimtime="00:00:31.87" resultid="12165" heatid="12741" lane="3" entrytime="00:00:31.04" entrycourse="SCM" />
                <RESULT eventid="1118" points="695" swimtime="00:05:59.23" resultid="12166" heatid="12769" lane="5" entrytime="00:06:20.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.17" />
                    <SPLIT distance="100" swimtime="00:01:20.50" />
                    <SPLIT distance="150" swimtime="00:02:10.32" />
                    <SPLIT distance="200" swimtime="00:02:58.06" />
                    <SPLIT distance="250" swimtime="00:03:47.19" />
                    <SPLIT distance="300" swimtime="00:04:37.89" />
                    <SPLIT distance="350" swimtime="00:05:19.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2190" points="652" swimtime="00:03:11.58" resultid="12167" heatid="12792" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.10" />
                    <SPLIT distance="100" swimtime="00:01:30.49" />
                    <SPLIT distance="150" swimtime="00:02:21.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CFP" nation="POR" region="ANNP" clubid="11991" name="Clube Fluvial Portuense" shortname="Fluvial Portuense">
          <ATHLETES>
            <ATHLETE firstname="Maria Fatima" lastname="Cabral" birthdate="1949-05-20" gender="F" nation="POR" license="106203" swrid="5048947" athleteid="12009">
              <RESULTS>
                <RESULT eventid="9659" status="DNS" swimtime="00:00:00.00" resultid="12010" heatid="12740" lane="8" entrytime="00:01:26.69" entrycourse="LCM" />
                <RESULT eventid="10350" status="DNS" swimtime="00:00:00.00" resultid="12011" heatid="12756" lane="2" entrytime="00:01:31.28" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Jorge" lastname="Marques" birthdate="1951-10-10" gender="M" nation="POR" license="130679" swrid="5001724" athleteid="12049">
              <RESULTS>
                <RESULT eventid="9685" points="231" swimtime="00:00:46.23" resultid="12050" heatid="12745" lane="3" entrytime="00:00:46.13" entrycourse="LCM" />
                <RESULT eventid="10364" points="228" swimtime="00:00:58.14" resultid="12051" heatid="12760" lane="1" entrytime="00:00:51.22" entrycourse="SCM" />
                <RESULT eventid="10426" points="221" swimtime="00:00:52.93" resultid="12052" heatid="12798" lane="4" entrytime="00:00:49.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabel Carolina" lastname="Neves" birthdate="1980-03-27" gender="F" nation="POR" license="202850" swrid="4889296" athleteid="12056">
              <RESULTS>
                <RESULT eventid="4102" points="327" swimtime="00:27:05.95" resultid="12057" heatid="12729" lane="4" entrytime="00:27:42.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.14" />
                    <SPLIT distance="100" swimtime="00:01:36.79" />
                    <SPLIT distance="150" swimtime="00:02:29.11" />
                    <SPLIT distance="200" swimtime="00:03:23.35" />
                    <SPLIT distance="250" swimtime="00:04:18.57" />
                    <SPLIT distance="300" swimtime="00:05:13.82" />
                    <SPLIT distance="350" swimtime="00:06:08.17" />
                    <SPLIT distance="400" swimtime="00:07:03.79" />
                    <SPLIT distance="450" swimtime="00:07:58.50" />
                    <SPLIT distance="500" swimtime="00:08:51.86" />
                    <SPLIT distance="550" swimtime="00:09:46.64" />
                    <SPLIT distance="600" swimtime="00:10:40.68" />
                    <SPLIT distance="650" swimtime="00:11:36.06" />
                    <SPLIT distance="700" swimtime="00:12:31.11" />
                    <SPLIT distance="750" swimtime="00:13:26.31" />
                    <SPLIT distance="800" swimtime="00:14:22.07" />
                    <SPLIT distance="850" swimtime="00:15:16.94" />
                    <SPLIT distance="900" swimtime="00:16:11.97" />
                    <SPLIT distance="950" swimtime="00:17:08.32" />
                    <SPLIT distance="1000" swimtime="00:18:03.14" />
                    <SPLIT distance="1050" swimtime="00:18:57.83" />
                    <SPLIT distance="1100" swimtime="00:19:52.44" />
                    <SPLIT distance="1150" swimtime="00:20:48.37" />
                    <SPLIT distance="1200" swimtime="00:21:47.16" />
                    <SPLIT distance="1250" swimtime="00:22:39.27" />
                    <SPLIT distance="1300" swimtime="00:23:35.01" />
                    <SPLIT distance="1400" swimtime="00:25:24.89" />
                    <SPLIT distance="1450" swimtime="00:26:18.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2111" points="241" swimtime="00:03:59.89" resultid="12058" heatid="12736" lane="2" entrytime="00:04:06.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.07" />
                    <SPLIT distance="100" swimtime="00:02:01.33" />
                    <SPLIT distance="150" swimtime="00:03:01.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2164" points="159" swimtime="00:01:59.05" resultid="12060" heatid="12750" lane="3" entrytime="00:01:54.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Miguel" lastname="Barroso" birthdate="1962-05-19" gender="M" nation="POR" license="208445" swrid="5326682" athleteid="11998">
              <RESULTS>
                <RESULT eventid="9685" points="706" swimtime="00:00:29.23" resultid="11999" heatid="12749" lane="5" entrytime="00:00:29.71" entrycourse="LCM" />
                <RESULT eventid="10364" points="591" swimtime="00:00:36.33" resultid="12000" heatid="12807" lane="7" entrytime="00:00:35.20" entrycourse="SCM" />
                <RESULT eventid="9789" points="630" swimtime="00:01:19.44" resultid="12001" heatid="12812" lane="3" entrytime="00:01:20.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Margarida Maria" lastname="Ribeiro" birthdate="1964-06-04" gender="F" nation="POR" license="131782" swrid="5036828" athleteid="12072">
              <RESULTS>
                <RESULT eventid="9659" points="180" swimtime="00:00:50.81" resultid="12073" heatid="12740" lane="3" entrytime="00:00:51.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos Guimaraes" lastname="Goncalves" birthdate="1970-11-22" gender="M" nation="POR" license="123664" swrid="4763854" athleteid="12037">
              <RESULTS>
                <RESULT eventid="2124" points="620" swimtime="00:02:43.15" resultid="12038" heatid="12737" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:20.14" />
                    <SPLIT distance="150" swimtime="00:02:01.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2177" points="688" swimtime="00:01:10.54" resultid="12039" heatid="12752" lane="2" entrytime="00:01:06.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="622" swimtime="00:05:52.59" resultid="12040" heatid="12770" lane="6" entrytime="00:05:45.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:14.36" />
                    <SPLIT distance="150" swimtime="00:02:00.43" />
                    <SPLIT distance="200" swimtime="00:02:46.22" />
                    <SPLIT distance="250" swimtime="00:03:38.42" />
                    <SPLIT distance="300" swimtime="00:04:32.32" />
                    <SPLIT distance="350" swimtime="00:05:13.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Goncalves" lastname="Costa" birthdate="1946-12-30" gender="M" nation="POR" license="131590" swrid="5030203" athleteid="12026">
              <RESULTS>
                <RESULT eventid="9685" points="184" swimtime="00:00:54.96" resultid="12027" heatid="12744" lane="4" entrytime="00:00:50.29" entrycourse="SCM" />
                <RESULT eventid="10364" points="205" swimtime="00:01:06.48" resultid="12028" heatid="12759" lane="3" entrytime="00:01:03.70" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Nuno" lastname="Goncalves" birthdate="1972-05-25" gender="M" nation="POR" license="205032" swrid="5227009" athleteid="12041">
              <RESULTS>
                <RESULT eventid="4128" status="DNS" swimtime="00:00:00.00" resultid="12042" heatid="12731" lane="8" entrytime="00:29:17.50" entrycourse="LCM" />
                <RESULT eventid="2177" status="DNS" swimtime="00:00:00.00" resultid="12043" heatid="12751" lane="6" entrytime="00:02:01.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Astride" lastname="Almeida" birthdate="1972-02-03" gender="F" nation="POR" license="212350" swrid="5424149" athleteid="11992">
              <RESULTS>
                <RESULT eventid="9711" status="DNS" swimtime="00:00:00.00" resultid="11993" heatid="12772" lane="2" entrytime="00:02:02.96" entrycourse="SCM" />
                <RESULT eventid="9763" status="DNS" swimtime="00:00:00.00" resultid="11994" heatid="12787" lane="6" entrytime="00:01:59.69" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ines Silva" lastname="Carvalho" birthdate="1983-08-16" gender="F" nation="POR" license="212606" swrid="5429040" athleteid="12016">
              <RESULTS>
                <RESULT eventid="2164" points="239" swimtime="00:01:42.65" resultid="12017" heatid="12750" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10350" points="306" swimtime="00:00:46.94" resultid="12018" heatid="12757" lane="6" entrytime="00:00:48.73" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elza Maria" lastname="Carvalho" birthdate="1976-01-13" gender="F" nation="POR" license="153144" swrid="5112926" athleteid="12012">
              <RESULTS>
                <RESULT eventid="9605" points="346" swimtime="00:01:36.60" resultid="12013" heatid="12804" lane="6" entrytime="00:01:33.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10350" points="489" swimtime="00:00:44.61" resultid="12014" heatid="12806" lane="8" entrytime="00:00:43.08" entrycourse="SCM" />
                <RESULT eventid="2190" points="517" swimtime="00:03:30.83" resultid="12015" heatid="12813" lane="6" entrytime="00:03:35.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.18" />
                    <SPLIT distance="100" swimtime="00:01:43.49" />
                    <SPLIT distance="150" swimtime="00:02:37.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Rui" lastname="Amaral" birthdate="1963-02-23" gender="M" nation="POR" license="206897" swrid="5276256" athleteid="11995">
              <RESULTS>
                <RESULT eventid="9685" status="DNS" swimtime="00:00:00.00" resultid="11996" heatid="12746" lane="5" entrytime="00:00:36.82" entrycourse="SCM" />
                <RESULT eventid="1157" points="332" swimtime="00:03:03.00" resultid="11997" heatid="12782" lane="7" entrytime="00:02:53.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.45" />
                    <SPLIT distance="100" swimtime="00:01:28.36" />
                    <SPLIT distance="150" swimtime="00:02:16.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Alves" lastname="Cecilio" birthdate="1954-04-10" gender="M" nation="POR" license="100919" swrid="4403439" athleteid="12022">
              <RESULTS>
                <RESULT eventid="9685" points="236" swimtime="00:00:44.58" resultid="12023" heatid="12745" lane="5" entrytime="00:00:42.43" entrycourse="SCM" />
                <RESULT eventid="10364" points="378" swimtime="00:00:46.93" resultid="12024" heatid="12762" lane="2" entrytime="00:00:42.60" entrycourse="SCM" />
                <RESULT eventid="10399" points="286" swimtime="00:00:50.54" resultid="12025" heatid="12786" lane="2" entrytime="00:00:48.41" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filipe Miguel" lastname="Silva" birthdate="1974-09-28" gender="M" nation="POR" license="201375" swrid="5171525" athleteid="12078">
              <RESULTS>
                <RESULT eventid="9632" points="193" swimtime="00:01:42.68" resultid="12079" heatid="12735" lane="3" entrytime="00:01:36.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.13" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="609 - O(A) nadador(a) não começou a executar a viragem imediatamente após terminar a braçada na posição ventral aos 50 metros - SW 6.4" eventid="2124" status="DSQ" swimtime="00:00:00.00" resultid="12080" heatid="12738" lane="1" entrytime="00:03:38.47" entrycourse="LCM" />
                <RESULT eventid="9685" points="289" swimtime="00:00:36.07" resultid="12081" heatid="12744" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Catarina Araujo" lastname="Blanco" birthdate="1971-11-08" gender="F" nation="POR" license="124701" swrid="4004822" athleteid="12005">
              <RESULTS>
                <RESULT eventid="9605" points="253" swimtime="00:01:46.18" resultid="12006" heatid="12804" lane="2" entrytime="00:01:36.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2111" points="281" swimtime="00:03:44.18" resultid="12007" heatid="12736" lane="5" entrytime="00:03:38.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.32" />
                    <SPLIT distance="100" swimtime="00:01:52.60" />
                    <SPLIT distance="150" swimtime="00:02:51.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10350" points="342" swimtime="00:00:51.17" resultid="12008" heatid="12757" lane="2" entrytime="00:00:49.08" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antero Silva" lastname="Sousa" birthdate="1943-10-16" gender="M" nation="POR" license="205243" swrid="5231633" athleteid="12082">
              <RESULTS>
                <RESULT eventid="9685" points="158" swimtime="00:00:57.83" resultid="12083" heatid="12744" lane="5" entrytime="00:00:56.25" entrycourse="LCM" />
                <RESULT eventid="10364" points="274" swimtime="00:01:00.35" resultid="12084" heatid="12759" lane="4" entrytime="00:00:55.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose Pedro" lastname="Neves" birthdate="1981-09-08" gender="M" nation="POR" license="17203" swrid="4190112" athleteid="12061">
              <RESULTS>
                <RESULT eventid="4128" status="DNS" swimtime="00:00:00.00" resultid="12062" heatid="12731" lane="5" entrytime="00:20:19.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Miguel" lastname="Bernardo" birthdate="1961-04-22" gender="M" nation="POR" license="201380" swrid="5171462" athleteid="12002">
              <RESULTS>
                <RESULT comment="Recorde Nacional " eventid="10364" points="697" swimtime="00:00:36.92" resultid="12003" heatid="12807" lane="8" entrytime="00:00:36.97" entrycourse="LCM" />
                <RESULT comment="Recorde Nacional " eventid="9789" points="688" swimtime="00:01:23.65" resultid="12004" heatid="12812" lane="2" entrytime="00:01:21.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo Francisco" lastname="Torres" birthdate="1962-11-12" gender="M" nation="POR" license="130665" swrid="5001750" athleteid="12087">
              <RESULTS>
                <RESULT eventid="4128" points="471" swimtime="00:22:36.41" resultid="12088" heatid="12731" lane="7" entrytime="00:23:36.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:22.31" />
                    <SPLIT distance="150" swimtime="00:02:06.90" />
                    <SPLIT distance="200" swimtime="00:02:51.43" />
                    <SPLIT distance="250" swimtime="00:03:36.47" />
                    <SPLIT distance="300" swimtime="00:04:21.46" />
                    <SPLIT distance="350" swimtime="00:05:06.89" />
                    <SPLIT distance="400" swimtime="00:05:52.00" />
                    <SPLIT distance="450" swimtime="00:06:37.23" />
                    <SPLIT distance="500" swimtime="00:07:22.27" />
                    <SPLIT distance="550" swimtime="00:08:08.03" />
                    <SPLIT distance="600" swimtime="00:08:52.90" />
                    <SPLIT distance="650" swimtime="00:09:38.74" />
                    <SPLIT distance="700" swimtime="00:10:23.54" />
                    <SPLIT distance="750" swimtime="00:11:09.63" />
                    <SPLIT distance="800" swimtime="00:11:54.44" />
                    <SPLIT distance="850" swimtime="00:12:40.11" />
                    <SPLIT distance="900" swimtime="00:13:25.99" />
                    <SPLIT distance="950" swimtime="00:14:11.69" />
                    <SPLIT distance="1000" swimtime="00:14:57.65" />
                    <SPLIT distance="1050" swimtime="00:15:43.00" />
                    <SPLIT distance="1100" swimtime="00:16:28.47" />
                    <SPLIT distance="1150" swimtime="00:17:16.30" />
                    <SPLIT distance="1200" swimtime="00:18:05.45" />
                    <SPLIT distance="1250" swimtime="00:18:50.41" />
                    <SPLIT distance="1300" swimtime="00:19:35.15" />
                    <SPLIT distance="1350" swimtime="00:20:21.13" />
                    <SPLIT distance="1400" swimtime="00:21:09.23" />
                    <SPLIT distance="1450" swimtime="00:21:52.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Miguel" lastname="Pinto" birthdate="1973-05-16" gender="M" nation="POR" license="208406" swrid="5326914" athleteid="12070">
              <RESULTS>
                <RESULT eventid="10364" points="349" swimtime="00:00:43.02" resultid="12071" heatid="12761" lane="3" entrytime="00:00:44.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Americo Pedro" lastname="Goncalves" birthdate="1971-05-19" gender="M" nation="POR" license="121758" swrid="4703094" athleteid="12034">
              <RESULTS>
                <RESULT eventid="2124" status="DNS" swimtime="00:00:00.00" resultid="12035" heatid="12738" lane="6" entrytime="00:02:36.68" entrycourse="SCM" />
                <RESULT eventid="9685" status="DNS" swimtime="00:00:00.00" resultid="12036" heatid="12805" lane="3" entrytime="00:00:26.62" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Alexandre" lastname="Inverneiro" birthdate="1971-04-21" gender="M" nation="POR" license="153118" swrid="5112952" athleteid="12044">
              <RESULTS>
                <RESULT eventid="9632" status="DNS" swimtime="00:00:00.00" resultid="12045" heatid="12735" lane="2" entrytime="00:01:42.16" entrycourse="SCM" />
                <RESULT eventid="2124" status="DNS" swimtime="00:00:00.00" resultid="12046" heatid="12738" lane="8" entrytime="00:03:45.76" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Maria" lastname="Cunha" birthdate="1971-09-03" gender="M" nation="POR" license="204079" swrid="4548183" athleteid="12031">
              <RESULTS>
                <RESULT eventid="9685" points="421" swimtime="00:00:32.98" resultid="12032" heatid="12748" lane="6" entrytime="00:00:33.11" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco David" lastname="Ferreira" birthdate="1989-07-25" gender="M" nation="POR" license="121874" swrid="4574825" athleteid="12033" />
            <ATHLETE firstname="Rui Alberto" lastname="Mendes" birthdate="1975-10-11" gender="M" nation="POR" license="202097" swrid="5197049" athleteid="12053">
              <RESULTS>
                <RESULT eventid="9632" points="296" swimtime="00:01:29.12" resultid="12054" heatid="12735" lane="4" entrytime="00:01:32.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9685" points="384" swimtime="00:00:32.84" resultid="12055" heatid="12748" lane="4" entrytime="00:00:32.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao Luis" lastname="Roseira" birthdate="1955-02-27" gender="M" nation="POR" license="142204" swrid="5119322" athleteid="12074">
              <RESULTS>
                <RESULT eventid="10364" points="149" swimtime="00:01:04.05" resultid="12075" heatid="12759" lane="5" entrytime="00:00:59.73" entrycourse="LCM" />
                <RESULT eventid="9737" points="143" swimtime="00:01:56.73" resultid="12076" heatid="12775" lane="2" entrytime="00:01:53.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="63" swimtime="00:01:16.42" resultid="12077" heatid="12798" lane="3" entrytime="00:01:04.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sergio Manuel" lastname="Neves" birthdate="1982-10-02" gender="M" nation="POR" license="204875" swrid="5215134" athleteid="12063">
              <RESULTS>
                <RESULT eventid="9737" points="195" swimtime="00:01:28.58" resultid="12064" heatid="12776" lane="2" entrytime="00:01:30.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="148" swimtime="00:03:30.35" resultid="12065" heatid="12781" lane="6" entrytime="00:03:39.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.27" />
                    <SPLIT distance="100" swimtime="00:01:42.14" />
                    <SPLIT distance="150" swimtime="00:02:37.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="114" swimtime="00:00:51.29" resultid="12066" heatid="12798" lane="5" entrytime="00:00:50.95" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nuno Silva" lastname="Lobo" birthdate="1963-12-13" gender="M" nation="POR" license="102544" swrid="5036815" athleteid="12047">
              <RESULTS>
                <RESULT eventid="9685" points="709" swimtime="00:00:29.18" resultid="12048" heatid="12749" lane="4" entrytime="00:00:28.63" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ivan Mauricio" lastname="Couras" birthdate="1981-02-08" gender="M" nation="POR" license="10232" swrid="4558833" athleteid="12029">
              <RESULTS>
                <RESULT eventid="4128" points="616" swimtime="00:19:31.56" resultid="12030" heatid="12731" lane="4" entrytime="00:19:16.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:12.63" />
                    <SPLIT distance="150" swimtime="00:01:50.67" />
                    <SPLIT distance="200" swimtime="00:02:28.81" />
                    <SPLIT distance="250" swimtime="00:03:06.87" />
                    <SPLIT distance="300" swimtime="00:03:45.12" />
                    <SPLIT distance="350" swimtime="00:04:23.73" />
                    <SPLIT distance="400" swimtime="00:05:02.52" />
                    <SPLIT distance="450" swimtime="00:05:41.31" />
                    <SPLIT distance="500" swimtime="00:06:19.75" />
                    <SPLIT distance="550" swimtime="00:06:58.45" />
                    <SPLIT distance="600" swimtime="00:07:37.32" />
                    <SPLIT distance="650" swimtime="00:08:16.13" />
                    <SPLIT distance="700" swimtime="00:08:55.11" />
                    <SPLIT distance="750" swimtime="00:09:34.18" />
                    <SPLIT distance="800" swimtime="00:10:13.79" />
                    <SPLIT distance="850" swimtime="00:10:53.68" />
                    <SPLIT distance="900" swimtime="00:11:33.30" />
                    <SPLIT distance="950" swimtime="00:12:13.09" />
                    <SPLIT distance="1000" swimtime="00:12:53.16" />
                    <SPLIT distance="1050" swimtime="00:13:33.10" />
                    <SPLIT distance="1100" swimtime="00:14:13.14" />
                    <SPLIT distance="1150" swimtime="00:14:53.15" />
                    <SPLIT distance="1200" swimtime="00:15:33.12" />
                    <SPLIT distance="1250" swimtime="00:16:13.30" />
                    <SPLIT distance="1300" swimtime="00:16:53.59" />
                    <SPLIT distance="1350" swimtime="00:17:33.76" />
                    <SPLIT distance="1400" swimtime="00:18:13.79" />
                    <SPLIT distance="1450" swimtime="00:18:53.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui David" lastname="Castro" birthdate="1970-04-03" gender="M" nation="POR" license="214263" swrid="5472931" athleteid="12019">
              <RESULTS>
                <RESULT eventid="9685" points="604" swimtime="00:00:29.23" resultid="12020" heatid="12805" lane="8" entrytime="00:00:29.15" entrycourse="LCM" />
                <RESULT eventid="2177" points="412" swimtime="00:01:23.68" resultid="12021" heatid="12752" lane="8" entrytime="00:01:16.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Abel" lastname="Pereira" birthdate="1973-11-12" gender="M" nation="POR" license="153155" swrid="5112981" athleteid="12067">
              <RESULTS>
                <RESULT eventid="9685" points="230" swimtime="00:00:38.93" resultid="12068" heatid="12746" lane="8" entrytime="00:00:42.07" entrycourse="SCM" />
                <RESULT eventid="2177" points="145" swimtime="00:01:51.25" resultid="12069" heatid="12751" lane="3" entrytime="00:01:46.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="10314" swimtime="00:02:41.94" resultid="12089" heatid="12803" lane="7" entrytime="00:02:38.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                    <SPLIT distance="100" swimtime="00:01:26.06" />
                    <SPLIT distance="150" swimtime="00:02:13.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12053" number="1" />
                    <RELAYPOSITION athleteid="12016" number="2" />
                    <RELAYPOSITION athleteid="12056" number="3" />
                    <RELAYPOSITION athleteid="12033" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="1061" swimtime="00:05:21.25" resultid="12090" heatid="12765" lane="6" entrytime="00:05:30.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:06.39" />
                    <SPLIT distance="150" swimtime="00:01:54.40" />
                    <SPLIT distance="200" swimtime="00:02:41.60" />
                    <SPLIT distance="250" swimtime="00:03:23.04" />
                    <SPLIT distance="300" swimtime="00:04:09.79" />
                    <SPLIT distance="350" swimtime="00:04:43.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12019" number="1" />
                    <RELAYPOSITION athleteid="12016" number="2" />
                    <RELAYPOSITION athleteid="12056" number="3" />
                    <RELAYPOSITION athleteid="12053" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="10378" status="DNS" swimtime="00:00:00.00" resultid="12091" heatid="12768" lane="6" entrytime="00:02:26.91">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11992" number="1" />
                    <RELAYPOSITION athleteid="11998" number="2" />
                    <RELAYPOSITION athleteid="12012" number="3" />
                    <RELAYPOSITION athleteid="12002" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="10314" swimtime="00:02:33.41" resultid="12092" heatid="12803" lane="4" entrytime="00:02:22.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                    <SPLIT distance="100" swimtime="00:01:22.51" />
                    <SPLIT distance="150" swimtime="00:01:54.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12029" number="1" />
                    <RELAYPOSITION athleteid="12012" number="2" />
                    <RELAYPOSITION athleteid="12037" number="3" />
                    <RELAYPOSITION athleteid="12005" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="2">
              <RESULTS>
                <RESULT eventid="1061" status="WDR" swimtime="00:00:00.00" resultid="12093" heatid="12765" lane="5" entrytime="00:04:40.15">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11998" number="1" />
                    <RELAYPOSITION athleteid="12005" number="2" />
                    <RELAYPOSITION athleteid="12012" number="3" />
                    <RELAYPOSITION athleteid="12034" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="319" agetotalmin="280" gender="X" number="3">
              <RESULTS>
                <RESULT eventid="10314" status="DNS" swimtime="00:00:00.00" resultid="12094" heatid="12728" lane="5" entrytime="00:04:24.38">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12082" number="1" />
                    <RELAYPOSITION athleteid="12009" number="2" />
                    <RELAYPOSITION athleteid="12072" number="3" />
                    <RELAYPOSITION athleteid="12026" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="CNPO" nation="POR" region="ANNP" clubid="11854" name="Clube Naval Povoense">
          <ATHLETES>
            <ATHLETE firstname="Marco Paulo" lastname="Silva" birthdate="1970-10-20" gender="M" nation="POR" license="118005" swrid="4577120" athleteid="11858">
              <RESULTS>
                <RESULT eventid="1157" points="324" swimtime="00:02:59.72" resultid="11859" heatid="12782" lane="2" entrytime="00:02:51.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                    <SPLIT distance="100" swimtime="00:01:23.91" />
                    <SPLIT distance="150" swimtime="00:02:13.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9789" points="355" swimtime="00:01:38.20" resultid="11860" heatid="12812" lane="8" entrytime="00:01:33.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Rosa" lastname="Serra" birthdate="1977-05-27" gender="F" nation="POR" license="205535" swrid="5260600" athleteid="11855">
              <RESULTS>
                <RESULT eventid="9711" points="163" swimtime="00:01:48.66" resultid="11856" heatid="12772" lane="3" entrytime="00:01:53.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9763" points="237" swimtime="00:02:02.27" resultid="11857" heatid="12787" lane="2" entrytime="00:02:06.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nuno Miguel" lastname="Silva" birthdate="1972-07-30" gender="M" nation="POR" license="206943" swrid="5277953" athleteid="11861">
              <RESULTS>
                <RESULT eventid="9737" points="283" swimtime="00:01:20.59" resultid="11862" heatid="12777" lane="8" entrytime="00:01:22.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="245" swimtime="00:03:03.33" resultid="11863" heatid="12781" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                    <SPLIT distance="100" swimtime="00:01:26.57" />
                    <SPLIT distance="150" swimtime="00:02:15.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CNMAL" nation="POR" region="ANL" clubid="11849" name="Clube Natacao Masters de Almada">
          <ATHLETES>
            <ATHLETE firstname="Ana Paula" lastname="Gonçalves" birthdate="1965-06-17" gender="F" nation="BRA" license="GB578407" swrid="5075614" athleteid="11850">
              <RESULTS>
                <RESULT eventid="2111" points="600" swimtime="00:03:15.00" resultid="11851" heatid="12736" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.38" />
                    <SPLIT distance="100" swimtime="00:01:34.27" />
                    <SPLIT distance="150" swimtime="00:02:25.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10386" points="536" swimtime="00:00:41.65" resultid="11852" heatid="12783" lane="7" />
                <RESULT eventid="10412" points="435" swimtime="00:00:42.14" resultid="11853" heatid="12795" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="FS" nation="POR" region="ANL" clubid="11877" name="Salesianos">
          <ATHLETES>
            <ATHLETE firstname="Alberto Vaz" lastname="Correia" birthdate="1955-09-22" gender="M" nation="POR" license="128374" swrid="4919450" athleteid="11878">
              <RESULTS>
                <RESULT comment="Recorde Nacional " eventid="4128" points="701" swimtime="00:22:36.53" resultid="11879" heatid="12731" lane="6" entrytime="00:22:41.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                    <SPLIT distance="100" swimtime="00:01:22.00" />
                    <SPLIT distance="150" swimtime="00:02:06.34" />
                    <SPLIT distance="200" swimtime="00:02:51.19" />
                    <SPLIT distance="250" swimtime="00:03:36.42" />
                    <SPLIT distance="300" swimtime="00:04:21.33" />
                    <SPLIT distance="350" swimtime="00:05:06.18" />
                    <SPLIT distance="400" swimtime="00:05:51.33" />
                    <SPLIT distance="450" swimtime="00:06:36.87" />
                    <SPLIT distance="500" swimtime="00:07:22.25" />
                    <SPLIT distance="550" swimtime="00:08:07.48" />
                    <SPLIT distance="600" swimtime="00:08:52.90" />
                    <SPLIT distance="650" swimtime="00:09:38.58" />
                    <SPLIT distance="700" swimtime="00:10:23.89" />
                    <SPLIT distance="750" swimtime="00:11:09.32" />
                    <SPLIT distance="800" swimtime="00:11:54.69" />
                    <SPLIT distance="850" swimtime="00:12:40.28" />
                    <SPLIT distance="900" swimtime="00:13:26.25" />
                    <SPLIT distance="950" swimtime="00:14:11.83" />
                    <SPLIT distance="1000" swimtime="00:14:57.67" />
                    <SPLIT distance="1050" swimtime="00:15:43.38" />
                    <SPLIT distance="1100" swimtime="00:16:29.29" />
                    <SPLIT distance="1150" swimtime="00:17:15.71" />
                    <SPLIT distance="1200" swimtime="00:18:02.26" />
                    <SPLIT distance="1250" swimtime="00:18:49.08" />
                    <SPLIT distance="1300" swimtime="00:19:35.50" />
                    <SPLIT distance="1350" swimtime="00:20:21.77" />
                    <SPLIT distance="1400" swimtime="00:21:08.03" />
                    <SPLIT distance="1450" swimtime="00:21:54.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9685" points="554" swimtime="00:00:33.58" resultid="11880" heatid="12748" lane="3" entrytime="00:00:31.44" entrycourse="SCM" />
                <RESULT eventid="1157" points="648" swimtime="00:02:44.89" resultid="11881" heatid="12782" lane="5" entrytime="00:02:36.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                    <SPLIT distance="100" swimtime="00:01:17.95" />
                    <SPLIT distance="150" swimtime="00:02:01.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="CNAL" nation="POR" region="ANDL" clubid="11928" name="Clube de Natacao de Alcobaca" shortname="Alcobaca">
          <ATHLETES>
            <ATHLETE firstname="Ana Rita" lastname="Freitas" birthdate="1986-12-26" gender="F" nation="POR" license="203951" swrid="5128536" athleteid="11933">
              <RESULTS>
                <RESULT eventid="9605" points="167" swimtime="00:01:59.56" resultid="11934" heatid="12733" lane="5" entrytime="00:01:54.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1144" points="204" swimtime="00:03:37.49" resultid="11935" heatid="12810" lane="1" entrytime="00:03:39.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.95" />
                    <SPLIT distance="100" swimtime="00:01:45.32" />
                    <SPLIT distance="150" swimtime="00:02:41.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10412" points="214" swimtime="00:00:47.54" resultid="11936" heatid="12795" lane="4" entrytime="00:00:49.86" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="David Jose" lastname="Oliveira" birthdate="1975-06-09" gender="M" nation="POR" license="203952" swrid="5128555" athleteid="11941">
              <RESULTS>
                <RESULT eventid="9632" points="117" swimtime="00:02:01.16" resultid="11942" heatid="12734" lane="4" entrytime="00:01:59.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9737" points="162" swimtime="00:01:37.00" resultid="11943" heatid="12775" lane="3" entrytime="00:01:37.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9789" points="119" swimtime="00:02:14.20" resultid="11944" heatid="12790" lane="2" entrytime="00:02:12.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel Filipe" lastname="Pimenta" birthdate="1995-02-23" gender="M" nation="POR" license="102300" swrid="4123939" athleteid="11945">
              <RESULTS>
                <RESULT eventid="9632" points="271" swimtime="00:01:25.00" resultid="11946" heatid="12734" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9737" points="247" swimtime="00:01:17.39" resultid="11947" heatid="12774" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9789" points="306" swimtime="00:01:31.97" resultid="11948" heatid="12789" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rui Marcal" lastname="Areias" birthdate="1975-01-17" gender="M" nation="POR" license="143386" swrid="5267469" athleteid="11929">
              <RESULTS>
                <RESULT eventid="9685" points="247" swimtime="00:00:38.00" resultid="11930" heatid="12746" lane="6" entrytime="00:00:38.06" entrycourse="SCM" />
                <RESULT eventid="10364" points="218" swimtime="00:00:50.32" resultid="11931" heatid="12761" lane="8" entrytime="00:00:48.56" entrycourse="SCM" />
                <RESULT eventid="2203" points="224" swimtime="00:04:02.88" resultid="11932" heatid="12794" lane="8" entrytime="00:03:45.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.43" />
                    <SPLIT distance="100" swimtime="00:01:55.87" />
                    <SPLIT distance="150" swimtime="00:02:58.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Patricia Sousa" lastname="Leal" birthdate="1977-03-18" gender="F" nation="POR" license="215231" athleteid="11937">
              <RESULTS>
                <RESULT eventid="9605" points="202" swimtime="00:01:55.72" resultid="11938" heatid="12733" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10350" points="279" swimtime="00:00:52.54" resultid="11939" heatid="12756" lane="8" />
                <RESULT eventid="9763" points="272" swimtime="00:01:56.70" resultid="11940" heatid="12787" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor Santos" lastname="Reis" birthdate="1970-02-13" gender="M" nation="POR" license="210274" swrid="5350246" athleteid="11949">
              <RESULTS>
                <RESULT eventid="9685" points="147" swimtime="00:00:46.74" resultid="11950" heatid="12745" lane="7" entrytime="00:00:49.54" entrycourse="SCM" />
                <RESULT eventid="10364" points="72" swimtime="00:01:13.66" resultid="11951" heatid="12758" lane="4" />
                <RESULT eventid="9737" points="110" swimtime="00:01:54.24" resultid="11952" heatid="12773" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="199" agetotalmin="160" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="10378" swimtime="00:02:53.91" resultid="11953" heatid="12767" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                    <SPLIT distance="100" swimtime="00:01:28.37" />
                    <SPLIT distance="150" swimtime="00:02:12.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11937" number="1" />
                    <RELAYPOSITION athleteid="11949" number="2" />
                    <RELAYPOSITION athleteid="11933" number="3" />
                    <RELAYPOSITION athleteid="11941" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="159" agetotalmin="120" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="10314" swimtime="00:03:00.79" resultid="11954" heatid="12728" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.80" />
                    <SPLIT distance="100" swimtime="00:01:44.07" />
                    <SPLIT distance="150" swimtime="00:02:19.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="11929" number="1" />
                    <RELAYPOSITION athleteid="11937" number="2" />
                    <RELAYPOSITION athleteid="11945" number="3" />
                    <RELAYPOSITION athleteid="11933" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="CNN" nation="POR" region="ANL" clubid="11955" name="Clube Nacional de Natação">
          <ATHLETES>
            <ATHLETE firstname="Paulo Gonçalves" lastname="Salvador" birthdate="1980-09-01" gender="M" nation="BRA" athleteid="11956">
              <RESULTS>
                <RESULT eventid="9685" points="599" swimtime="00:00:27.52" resultid="11957" heatid="12742" lane="4" />
                <RESULT eventid="9737" points="610" swimtime="00:01:00.44" resultid="11958" heatid="12773" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="535" swimtime="00:02:19.18" resultid="11959" heatid="12779" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                    <SPLIT distance="100" swimtime="00:01:06.98" />
                    <SPLIT distance="150" swimtime="00:01:44.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="FOCA" nation="POR" region="ANNP" clubid="12095" name="Foca-Clube de Natação de Felgueiras" shortname="Foca">
          <ATHLETES>
            <ATHLETE firstname="Vitorino Fernando" lastname="Faria" birthdate="1973-01-01" gender="M" nation="POR" license="147080" swrid="5091481" athleteid="12100">
              <RESULTS>
                <RESULT eventid="1157" points="186" swimtime="00:03:20.83" resultid="12101" heatid="12781" lane="4" entrytime="00:03:14.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.75" />
                    <SPLIT distance="100" swimtime="00:01:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="183" swimtime="00:00:45.21" resultid="12102" heatid="12799" lane="2" entrytime="00:00:44.54" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Rosa" lastname="Silva" birthdate="1980-11-19" gender="F" nation="POR" license="133361" swrid="5087251" athleteid="12128">
              <RESULTS>
                <RESULT eventid="2111" points="239" swimtime="00:04:00.41" resultid="12129" heatid="12736" lane="6" entrytime="00:03:56.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.92" />
                    <SPLIT distance="100" swimtime="00:01:57.63" />
                    <SPLIT distance="150" swimtime="00:02:59.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1118" points="672" swimtime="00:06:03.36" resultid="12130" heatid="12769" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.66" />
                    <SPLIT distance="100" swimtime="00:01:51.04" />
                    <SPLIT distance="200" swimtime="00:03:54.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rosa Leitao" lastname="Costa" birthdate="1965-07-15" gender="F" nation="POR" license="132419" swrid="5068113" athleteid="12096">
              <RESULTS>
                <RESULT eventid="9659" points="157" swimtime="00:00:53.19" resultid="12097" heatid="12740" lane="2" entrytime="00:00:54.64" entrycourse="LCM" />
                <RESULT eventid="10350" points="290" swimtime="00:00:56.71" resultid="12098" heatid="12756" lane="3" entrytime="00:00:54.77" entrycourse="SCM" />
                <RESULT eventid="2190" points="393" swimtime="00:04:12.88" resultid="12099" heatid="12813" lane="7" entrytime="00:04:01.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.40" />
                    <SPLIT distance="100" swimtime="00:02:01.34" />
                    <SPLIT distance="150" swimtime="00:03:07.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor Carvalho" lastname="Lopes" birthdate="1972-09-24" gender="M" nation="POR" license="132421" swrid="5068135" athleteid="12109">
              <RESULTS>
                <RESULT eventid="9737" status="DNS" swimtime="00:00:00.00" resultid="12110" heatid="12776" lane="7" entrytime="00:01:31.37" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Manuel" lastname="Ribeiro" birthdate="1991-07-27" gender="M" nation="POR" license="107830" swrid="5326937" athleteid="12121">
              <RESULTS>
                <RESULT eventid="9685" points="514" swimtime="00:00:27.61" resultid="12122" heatid="12805" lane="6" entrytime="00:00:28.01" entrycourse="LCM" />
                <RESULT eventid="1157" points="448" swimtime="00:02:19.11" resultid="12123" heatid="12811" lane="3" entrytime="00:02:27.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:06.23" />
                    <SPLIT distance="150" swimtime="00:01:43.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="402" swimtime="00:00:30.97" resultid="12124" heatid="12800" lane="5" entrytime="00:00:33.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuel Fernando" lastname="Fernandes" birthdate="1968-03-14" gender="M" nation="POR" license="202748" swrid="4845987" athleteid="12103">
              <RESULTS>
                <RESULT eventid="9685" points="115" swimtime="00:00:50.70" resultid="12104" heatid="12745" lane="8" entrytime="00:00:49.77" entrycourse="SCM" />
                <RESULT eventid="10364" points="188" swimtime="00:00:53.64" resultid="12105" heatid="12760" lane="7" entrytime="00:00:52.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Cunha" lastname="Ribeiro" birthdate="1970-01-22" gender="M" nation="POR" license="153289" swrid="5115801" athleteid="12125">
              <RESULTS>
                <RESULT eventid="9737" points="202" swimtime="00:01:33.18" resultid="12126" heatid="12776" lane="6" entrytime="00:01:30.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="262" swimtime="00:00:42.74" resultid="12127" heatid="12799" lane="7" entrytime="00:00:44.58" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filipe Pinheiro" lastname="Pires" birthdate="1973-05-02" gender="M" nation="POR" license="117638" swrid="4557827" athleteid="12119">
              <RESULTS>
                <RESULT eventid="2124" points="395" swimtime="00:02:59.30" resultid="12120" heatid="12738" lane="2" entrytime="00:02:46.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.36" />
                    <SPLIT distance="100" swimtime="00:01:29.49" />
                    <SPLIT distance="150" swimtime="00:02:15.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Filipe" lastname="Pimentel" birthdate="1984-01-22" gender="M" nation="POR" license="101691" swrid="5068153" athleteid="12117">
              <RESULTS>
                <RESULT eventid="1131" points="493" swimtime="00:05:45.43" resultid="12118" heatid="12770" lane="5" entrytime="00:05:34.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:14.10" />
                    <SPLIT distance="150" swimtime="00:01:59.08" />
                    <SPLIT distance="200" swimtime="00:02:41.79" />
                    <SPLIT distance="250" swimtime="00:03:31.43" />
                    <SPLIT distance="300" swimtime="00:04:20.87" />
                    <SPLIT distance="350" swimtime="00:05:03.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mario Nuno" lastname="Pereira" birthdate="1981-02-20" gender="M" nation="POR" license="200652" swrid="5157491" athleteid="12114">
              <RESULTS>
                <RESULT eventid="1157" points="336" swimtime="00:02:42.43" resultid="12115" heatid="12811" lane="8" entrytime="00:02:34.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                    <SPLIT distance="100" swimtime="00:01:13.89" />
                    <SPLIT distance="150" swimtime="00:01:58.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="411" swimtime="00:00:33.79" resultid="12116" heatid="12800" lane="3" entrytime="00:00:33.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose" lastname="Leite" birthdate="1948-09-16" gender="M" nation="POR" license="204547" swrid="5207388" athleteid="12106">
              <RESULTS>
                <RESULT eventid="9685" points="201" swimtime="00:00:48.45" resultid="12107" heatid="12745" lane="2" entrytime="00:00:45.45" entrycourse="SCM" />
                <RESULT eventid="2203" points="362" swimtime="00:04:19.83" resultid="12108" heatid="12793" lane="5" entrytime="00:04:18.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.01" />
                    <SPLIT distance="100" swimtime="00:02:05.30" />
                    <SPLIT distance="150" swimtime="00:03:14.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Catarina" lastname="Teixeira" birthdate="1995-02-16" gender="F" nation="POR" license="18137" swrid="4123386" athleteid="12135">
              <RESULTS>
                <RESULT eventid="9659" points="469" swimtime="00:00:32.54" resultid="12136" heatid="12741" lane="2" entrytime="00:00:33.01" entrycourse="SCM" />
                <RESULT eventid="10350" points="430" swimtime="00:00:41.84" resultid="12137" heatid="12755" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Albano Couto" lastname="Teixeira" birthdate="1963-08-30" gender="M" nation="POR" license="117114" swrid="5068174" athleteid="12131">
              <RESULTS>
                <RESULT eventid="9685" points="181" swimtime="00:00:45.96" resultid="12132" heatid="12745" lane="1" entrytime="00:00:49.73" entrycourse="SCM" />
                <RESULT eventid="10364" points="196" swimtime="00:00:52.49" resultid="12133" heatid="12760" lane="6" entrytime="00:00:50.06" entrycourse="SCM" />
                <RESULT eventid="2203" points="227" swimtime="00:04:25.54" resultid="12134" heatid="12793" lane="3" entrytime="00:04:20.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.15" />
                    <SPLIT distance="100" swimtime="00:02:06.26" />
                    <SPLIT distance="150" swimtime="00:03:17.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro Filipe" lastname="Martins" birthdate="1990-11-12" gender="M" nation="POR" license="22442" swrid="4559626" athleteid="12111">
              <RESULTS>
                <RESULT eventid="1157" points="498" swimtime="00:02:14.36" resultid="12112" heatid="12781" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.32" />
                    <SPLIT distance="100" swimtime="00:01:03.33" />
                    <SPLIT distance="150" swimtime="00:01:38.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="384" swimtime="00:00:31.45" resultid="12113" heatid="12797" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="SCE" nation="POR" region="ANCNP" clubid="12559" name="Sporting Clube de Espinho" shortname="Sporting de Espinho">
          <ATHLETES>
            <ATHLETE firstname="Maria Manuela" lastname="Oliveira" birthdate="1974-11-07" gender="F" nation="POR" license="208451" swrid="5326883" athleteid="12576">
              <RESULTS>
                <RESULT eventid="2111" points="324" swimtime="00:03:43.83" resultid="12701" heatid="12736" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.78" />
                    <SPLIT distance="100" swimtime="00:01:48.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10350" points="330" swimtime="00:00:50.88" resultid="12702" heatid="12757" lane="3" entrytime="00:00:48.05" entrycourse="SCM" />
                <RESULT eventid="9711" points="284" swimtime="00:01:30.66" resultid="12703" heatid="12808" lane="2" entrytime="00:01:27.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabio" lastname="Floriano" birthdate="1963-10-07" gender="M" nation="POR" license="207665" swrid="5297527" athleteid="12572">
              <RESULTS>
                <RESULT eventid="9685" points="339" swimtime="00:00:37.32" resultid="12573" heatid="12747" lane="1" entrytime="00:00:34.62" entrycourse="SCM" />
                <RESULT eventid="10364" points="301" swimtime="00:00:45.50" resultid="12574" heatid="12762" lane="1" entrytime="00:00:43.29" entrycourse="SCM" />
                <RESULT eventid="1157" points="263" swimtime="00:03:17.72" resultid="12575" heatid="12781" lane="5" entrytime="00:03:16.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                    <SPLIT distance="100" swimtime="00:01:30.72" />
                    <SPLIT distance="150" swimtime="00:02:25.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Domingos Jose" lastname="Ferreira" birthdate="1954-11-05" gender="M" nation="POR" license="209351" swrid="5336707" athleteid="12568">
              <RESULTS>
                <RESULT eventid="9737" points="305" swimtime="00:01:30.75" resultid="12569" heatid="12776" lane="4" entrytime="00:01:27.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="364" swimtime="00:03:19.78" resultid="12570" heatid="12782" lane="8" entrytime="00:03:13.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.27" />
                    <SPLIT distance="100" swimtime="00:01:33.30" />
                    <SPLIT distance="150" swimtime="00:02:26.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2203" points="391" swimtime="00:04:08.47" resultid="12571" heatid="12793" lane="4" entrytime="00:03:59.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.09" />
                    <SPLIT distance="100" swimtime="00:02:00.17" />
                    <SPLIT distance="150" swimtime="00:03:04.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yolanda" lastname="Rienderhoff" birthdate="1979-07-04" gender="F" nation="POR" license="207733" swrid="4886320" athleteid="12577">
              <RESULTS>
                <RESULT eventid="9659" status="DNS" swimtime="00:00:00.00" resultid="12578" heatid="12741" lane="7" entrytime="00:00:34.90" entrycourse="LCM" />
                <RESULT eventid="9711" points="410" swimtime="00:01:19.94" resultid="12579" heatid="12808" lane="4" entrytime="00:01:16.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2190" points="455" swimtime="00:03:35.95" resultid="12580" heatid="12813" lane="3" entrytime="00:03:28.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.92" />
                    <SPLIT distance="100" swimtime="00:01:43.31" />
                    <SPLIT distance="150" swimtime="00:02:41.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis Alberto" lastname="Esparragoza" birthdate="1980-04-19" gender="M" nation="POR" license="213246" swrid="5448493" athleteid="12564">
              <RESULTS>
                <RESULT eventid="9685" points="406" swimtime="00:00:31.34" resultid="12565" heatid="12749" lane="8" entrytime="00:00:31.06" entrycourse="SCM" />
                <RESULT eventid="10364" points="374" swimtime="00:00:40.36" resultid="12566" heatid="12759" lane="8" />
                <RESULT eventid="1157" points="390" swimtime="00:02:34.66" resultid="12567" heatid="12780" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                    <SPLIT distance="100" swimtime="00:01:14.15" />
                    <SPLIT distance="150" swimtime="00:01:55.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio Monteiro" lastname="Canelas" birthdate="1950-01-26" gender="M" nation="POR" license="148547" swrid="5100108" athleteid="12560">
              <RESULTS>
                <RESULT eventid="9737" points="244" swimtime="00:01:43.36" resultid="12561" heatid="12775" lane="4" entrytime="00:01:40.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9789" points="333" swimtime="00:01:58.94" resultid="12562" heatid="12790" lane="4" entrytime="00:01:50.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10426" points="262" swimtime="00:00:50.04" resultid="12563" heatid="12799" lane="1" entrytime="00:00:44.70" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuel Rui" lastname="Sousa" birthdate="1980-09-21" gender="M" nation="POR" license="213247" swrid="5448494" athleteid="12581">
              <RESULTS>
                <RESULT eventid="9685" points="256" swimtime="00:00:36.54" resultid="12582" heatid="12744" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="239" agetotalmin="200" gender="X" number="1">
              <RESULTS>
                <RESULT eventid="10378" swimtime="00:02:39.29" resultid="12583" heatid="12768" lane="2" entrytime="00:02:27.93">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                    <SPLIT distance="100" swimtime="00:01:23.75" />
                    <SPLIT distance="150" swimtime="00:01:58.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="12576" number="1" />
                    <RELAYPOSITION athleteid="12560" number="2" />
                    <RELAYPOSITION athleteid="12577" number="3" />
                    <RELAYPOSITION athleteid="12568" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="CCLV" nation="POR" region="ANL" clubid="11764" name="Clube de Campismo Luz e Vida">
          <ATHLETES>
            <ATHLETE firstname="Mário Nuno" lastname="Lopes" birthdate="1974-09-28" gender="M" nation="POR" license="212131" athleteid="11772">
              <RESULTS>
                <RESULT eventid="9632" status="DNS" swimtime="00:00:00.00" resultid="11773" heatid="12734" lane="7" />
                <RESULT eventid="9737" status="DNS" swimtime="00:00:00.00" resultid="11774" heatid="12773" lane="8" />
                <RESULT eventid="10426" status="DNS" swimtime="00:00:00.00" resultid="11775" heatid="12797" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana Filipa" lastname="Prior" birthdate="1977-08-29" gender="F" nation="POR" license="105895" swrid="5326294" athleteid="11765">
              <RESULTS>
                <RESULT eventid="4102" status="DNS" swimtime="00:00:00.00" resultid="11766" heatid="12729" lane="3" />
                <RESULT eventid="2111" status="DNS" swimtime="00:00:00.00" resultid="11767" heatid="12736" lane="4" entrytime="00:02:59.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno Gonçalo" lastname="Campos" birthdate="1976-11-12" gender="M" nation="POR" license="206910" swrid="5276195" athleteid="11768">
              <RESULTS>
                <RESULT eventid="9685" status="DNS" swimtime="00:00:00.00" resultid="11769" heatid="12748" lane="2" entrytime="00:00:33.28" entrycourse="LCM" />
                <RESULT eventid="10364" status="DNS" swimtime="00:00:00.00" resultid="11770" heatid="12763" lane="1" entrytime="00:00:41.96" entrycourse="SCM" />
                <RESULT eventid="10399" status="DNS" swimtime="00:00:00.00" resultid="11771" heatid="12786" lane="3" entrytime="00:00:42.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="VSC" nation="POR" region="ANNP" clubid="12598" name="Vitória Sport Clube">
          <ATHLETES>
            <ATHLETE firstname="Jose Orlando" lastname="Novais" birthdate="1978-10-20" gender="M" nation="POR" license="110370" swrid="4372968" athleteid="12610">
              <RESULTS>
                <RESULT eventid="9685" points="278" swimtime="00:00:35.56" resultid="12611" heatid="12747" lane="2" entrytime="00:00:34.36" entrycourse="SCM" />
                <RESULT eventid="9737" points="259" swimtime="00:01:20.41" resultid="12612" heatid="12773" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9789" points="316" swimtime="00:01:33.35" resultid="12613" heatid="12812" lane="1" entrytime="00:01:31.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Norberto Matos" lastname="Pereira" birthdate="1975-10-18" gender="M" nation="POR" license="111733" swrid="4403592" athleteid="12614">
              <RESULTS>
                <RESULT eventid="9737" status="WDR" swimtime="00:00:00.00" resultid="12615" heatid="12777" lane="3" entrytime="00:01:20.73" entrycourse="LCM" />
                <RESULT eventid="9789" status="WDR" swimtime="00:00:00.00" resultid="12616" heatid="12790" lane="3" entrytime="00:01:51.25" entrycourse="SCM" />
                <RESULT eventid="10426" status="WDR" swimtime="00:00:00.00" resultid="12617" heatid="12799" lane="8" entrytime="00:00:49.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agostinho Jorge" lastname="Sousa" birthdate="1981-09-21" gender="M" nation="POR" license="203962" swrid="5125755" athleteid="12618">
              <RESULTS>
                <RESULT eventid="9685" points="236" swimtime="00:00:37.52" resultid="12619" heatid="12747" lane="5" entrytime="00:00:35.22" entrycourse="LCM" />
                <RESULT eventid="10364" points="255" swimtime="00:00:45.82" resultid="12620" heatid="12761" lane="6" entrytime="00:00:46.10" entrycourse="LCM" />
                <RESULT eventid="9737" points="156" swimtime="00:01:35.21" resultid="12621" heatid="12776" lane="1" entrytime="00:01:32.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria Manuela" lastname="Ferreira" birthdate="1970-07-16" gender="F" nation="POR" license="130114" swrid="4988912" athleteid="12599">
              <RESULTS>
                <RESULT eventid="10322" points="134" swimtime="00:04:53.39" resultid="12600" heatid="12753" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.19" />
                    <SPLIT distance="100" swimtime="00:02:13.21" />
                    <SPLIT distance="150" swimtime="00:03:32.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="9711" points="317" swimtime="00:01:29.29" resultid="12601" heatid="12808" lane="7" entrytime="00:01:28.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="10412" points="195" swimtime="00:00:53.65" resultid="12602" heatid="12795" lane="5" entrytime="00:00:51.73" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Armindo Manuel" lastname="Lobo" birthdate="1984-04-17" gender="M" nation="POR" license="118906" swrid="4590317" athleteid="12606">
              <RESULTS>
                <RESULT eventid="9685" status="WDR" swimtime="00:00:00.00" resultid="12607" heatid="12805" lane="1" entrytime="00:00:29.13" entrycourse="LCM" />
                <RESULT eventid="9737" status="WDR" swimtime="00:00:00.00" resultid="12608" heatid="12809" lane="6" entrytime="00:01:02.82" entrycourse="SCM" />
                <RESULT eventid="10426" status="WDR" swimtime="00:00:00.00" resultid="12609" heatid="12800" lane="4" entrytime="00:00:31.77" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edgar Manuel" lastname="Guimaraes" birthdate="1980-09-10" gender="M" nation="POR" license="110317" swrid="4372958" athleteid="12603">
              <RESULTS>
                <RESULT eventid="9685" points="307" swimtime="00:00:34.40" resultid="12604" heatid="12748" lane="7" entrytime="00:00:33.28" entrycourse="LCM" />
                <RESULT eventid="10364" points="339" swimtime="00:00:41.68" resultid="12605" heatid="12763" lane="6" entrytime="00:00:40.94" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
  <TIMESTANDARDLISTS>
    <TIMESTANDARDLIST timestandardlistid="10455" code="01" course="SCM" gender="F" name="Masters FEM" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="25" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:27:30.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="10441" code="01" course="SCM" gender="M" name="Masters Masc" type="MAXIMUM">
      <AGEGROUP agemax="-1" agemin="25" />
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:25:00.00">
          <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:00.00">
          <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
  </TIMESTANDARDLISTS>
</LENEX>
